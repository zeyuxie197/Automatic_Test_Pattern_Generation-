1 1 0 2 0
2 13 1 1
2 14 1 1
1 4 0 2 0
2 15 1 4
2 16 1 4
1 7 0 2 0
2 17 1 7
2 18 1 7
1 10 0 2 0
2 19 1 10
2 20 1 10
0 21 5 1 1 13
0 22 7 2 2 16 17
2 26 1 22
2 27 1 22
0 25 5 1 1 20
0 28 6 1 2 15 21
0 29 6 1 2 14 26
0 30 6 1 2 27 19
0 31 6 1 2 25 18
3 32 6 0 4 28 29 30 31