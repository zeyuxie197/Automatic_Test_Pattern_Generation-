1 1 0 16 0 
2 2 1 1  
2 3 1 1  
2 4 1 1  
2 5 1 1  
2 6 1 1  
2 7 1 1  
2 8 1 1  
2 9 1 1  
2 10 1 1  
2 11 1 1  
2 12 1 1  
2 13 1 1  
2 14 1 1  
2 15 1 1  
2 16 1 1  
2 17 1 1  
1 18 0 16 0 
2 19 1 18  
2 20 1 18  
2 21 1 18  
2 22 1 18  
2 23 1 18  
2 24 1 18  
2 25 1 18  
2 26 1 18  
2 27 1 18  
2 28 1 18  
2 29 1 18  
2 30 1 18  
2 31 1 18  
2 32 1 18  
2 33 1 18  
2 34 1 18  
1 35 0 16 0 
2 36 1 35  
2 37 1 35  
2 38 1 35  
2 39 1 35  
2 40 1 35  
2 41 1 35  
2 42 1 35  
2 43 1 35  
2 44 1 35  
2 45 1 35  
2 46 1 35  
2 47 1 35  
2 48 1 35  
2 49 1 35  
2 50 1 35  
2 51 1 35  
1 52 0 16 0 
2 53 1 52  
2 54 1 52  
2 55 1 52  
2 56 1 52  
2 57 1 52  
2 58 1 52  
2 59 1 52  
2 60 1 52  
2 61 1 52  
2 62 1 52  
2 63 1 52  
2 64 1 52  
2 65 1 52  
2 66 1 52  
2 67 1 52  
2 68 1 52  
1 69 0 16 0 
2 70 1 69  
2 71 1 69  
2 72 1 69  
2 73 1 69  
2 74 1 69  
2 75 1 69  
2 76 1 69  
2 77 1 69  
2 78 1 69  
2 79 1 69  
2 80 1 69  
2 81 1 69  
2 82 1 69  
2 83 1 69  
2 84 1 69  
2 85 1 69  
1 86 0 16 0 
2 87 1 86  
2 88 1 86  
2 89 1 86  
2 90 1 86  
2 91 1 86  
2 92 1 86  
2 93 1 86  
2 94 1 86  
2 95 1 86  
2 96 1 86  
2 97 1 86  
2 98 1 86  
2 99 1 86  
2 100 1 86  
2 101 1 86  
2 102 1 86  
1 103 0 16 0 
2 104 1 103  
2 105 1 103  
2 106 1 103  
2 107 1 103  
2 108 1 103  
2 109 1 103  
2 110 1 103  
2 111 1 103  
2 112 1 103  
2 113 1 103  
2 114 1 103  
2 115 1 103  
2 116 1 103  
2 117 1 103  
2 118 1 103  
2 119 1 103  
1 120 0 16 0 
2 121 1 120  
2 122 1 120  
2 123 1 120  
2 124 1 120  
2 125 1 120  
2 126 1 120  
2 127 1 120  
2 128 1 120  
2 129 1 120  
2 130 1 120  
2 131 1 120  
2 132 1 120  
2 133 1 120  
2 134 1 120  
2 135 1 120  
2 136 1 120  
1 137 0 16 0 
2 138 1 137  
2 139 1 137  
2 140 1 137  
2 141 1 137  
2 142 1 137  
2 143 1 137  
2 144 1 137  
2 145 1 137  
2 146 1 137  
2 147 1 137  
2 148 1 137  
2 149 1 137  
2 150 1 137  
2 151 1 137  
2 152 1 137  
2 153 1 137  
1 154 0 16 0 
2 155 1 154  
2 156 1 154  
2 157 1 154  
2 158 1 154  
2 159 1 154  
2 160 1 154  
2 161 1 154  
2 162 1 154  
2 163 1 154  
2 164 1 154  
2 165 1 154  
2 166 1 154  
2 167 1 154  
2 168 1 154  
2 169 1 154  
2 170 1 154  
1 171 0 16 0 
2 172 1 171  
2 173 1 171  
2 174 1 171  
2 175 1 171  
2 176 1 171  
2 177 1 171  
2 178 1 171  
2 179 1 171  
2 180 1 171  
2 181 1 171  
2 182 1 171  
2 183 1 171  
2 184 1 171  
2 185 1 171  
2 186 1 171  
2 187 1 171  
1 188 0 16 0 
2 189 1 188  
2 190 1 188  
2 191 1 188  
2 192 1 188  
2 193 1 188  
2 194 1 188  
2 195 1 188  
2 196 1 188  
2 197 1 188  
2 198 1 188  
2 199 1 188  
2 200 1 188  
2 201 1 188  
2 202 1 188  
2 203 1 188  
2 204 1 188  
1 205 0 16 0 
2 206 1 205  
2 207 1 205  
2 208 1 205  
2 209 1 205  
2 210 1 205  
2 211 1 205  
2 212 1 205  
2 213 1 205  
2 214 1 205  
2 215 1 205  
2 216 1 205  
2 217 1 205  
2 218 1 205  
2 219 1 205  
2 220 1 205  
2 221 1 205  
1 222 0 16 0 
2 223 1 222  
2 224 1 222  
2 225 1 222  
2 226 1 222  
2 227 1 222  
2 228 1 222  
2 229 1 222  
2 230 1 222  
2 231 1 222  
2 232 1 222  
2 233 1 222  
2 234 1 222  
2 235 1 222  
2 236 1 222  
2 237 1 222  
2 238 1 222  
1 239 0 16 0 
2 240 1 239  
2 241 1 239  
2 242 1 239  
2 243 1 239  
2 244 1 239  
2 245 1 239  
2 246 1 239  
2 247 1 239  
2 248 1 239  
2 249 1 239  
2 250 1 239  
2 251 1 239  
2 252 1 239  
2 253 1 239  
2 254 1 239  
2 255 1 239  
1 256 0 16 0 
2 257 1 256  
2 258 1 256  
2 259 1 256  
2 260 1 256  
2 261 1 256  
2 262 1 256  
2 263 1 256  
2 264 1 256  
2 265 1 256  
2 266 1 256  
2 267 1 256  
2 268 1 256  
2 269 1 256  
2 270 1 256  
2 271 1 256  
2 272 1 256  
1 273 0 16 0 
2 274 1 273  
2 275 1 273  
2 276 1 273  
2 277 1 273  
2 278 1 273  
2 279 1 273  
2 280 1 273  
2 281 1 273  
2 282 1 273  
2 283 1 273  
2 284 1 273  
2 285 1 273  
2 286 1 273  
2 287 1 273  
2 288 1 273  
2 289 1 273  
1 290 0 16 0 
2 291 1 290  
2 292 1 290  
2 293 1 290  
2 294 1 290  
2 295 1 290  
2 296 1 290  
2 297 1 290  
2 298 1 290  
2 299 1 290  
2 300 1 290  
2 301 1 290  
2 302 1 290  
2 303 1 290  
2 304 1 290  
2 305 1 290  
2 306 1 290  
1 307 0 16 0 
2 308 1 307  
2 309 1 307  
2 310 1 307  
2 311 1 307  
2 312 1 307  
2 313 1 307  
2 314 1 307  
2 315 1 307  
2 316 1 307  
2 317 1 307  
2 318 1 307  
2 319 1 307  
2 320 1 307  
2 321 1 307  
2 322 1 307  
2 323 1 307  
1 324 0 16 0 
2 325 1 324  
2 326 1 324  
2 327 1 324  
2 328 1 324  
2 329 1 324  
2 330 1 324  
2 331 1 324  
2 332 1 324  
2 333 1 324  
2 334 1 324  
2 335 1 324  
2 336 1 324  
2 337 1 324  
2 338 1 324  
2 339 1 324  
2 340 1 324  
1 341 0 16 0 
2 342 1 341  
2 343 1 341  
2 344 1 341  
2 345 1 341  
2 346 1 341  
2 347 1 341  
2 348 1 341  
2 349 1 341  
2 350 1 341  
2 351 1 341  
2 352 1 341  
2 353 1 341  
2 354 1 341  
2 355 1 341  
2 356 1 341  
2 357 1 341  
1 358 0 16 0 
2 359 1 358  
2 360 1 358  
2 361 1 358  
2 362 1 358  
2 363 1 358  
2 364 1 358  
2 365 1 358  
2 366 1 358  
2 367 1 358  
2 368 1 358  
2 369 1 358  
2 370 1 358  
2 371 1 358  
2 372 1 358  
2 373 1 358  
2 374 1 358  
1 375 0 16 0 
2 376 1 375  
2 377 1 375  
2 378 1 375  
2 379 1 375  
2 380 1 375  
2 381 1 375  
2 382 1 375  
2 383 1 375  
2 384 1 375  
2 385 1 375  
2 386 1 375  
2 387 1 375  
2 388 1 375  
2 389 1 375  
2 390 1 375  
2 391 1 375  
1 392 0 16 0 
2 393 1 392  
2 394 1 392  
2 395 1 392  
2 396 1 392  
2 397 1 392  
2 398 1 392  
2 399 1 392  
2 400 1 392  
2 401 1 392  
2 402 1 392  
2 403 1 392  
2 404 1 392  
2 405 1 392  
2 406 1 392  
2 407 1 392  
2 408 1 392  
1 409 0 16 0 
2 410 1 409  
2 411 1 409  
2 412 1 409  
2 413 1 409  
2 414 1 409  
2 415 1 409  
2 416 1 409  
2 417 1 409  
2 418 1 409  
2 419 1 409  
2 420 1 409  
2 421 1 409  
2 422 1 409  
2 423 1 409  
2 424 1 409  
2 425 1 409  
1 426 0 16 0 
2 427 1 426  
2 428 1 426  
2 429 1 426  
2 430 1 426  
2 431 1 426  
2 432 1 426  
2 433 1 426  
2 434 1 426  
2 435 1 426  
2 436 1 426  
2 437 1 426  
2 438 1 426  
2 439 1 426  
2 440 1 426  
2 441 1 426  
2 442 1 426  
1 443 0 16 0 
2 444 1 443  
2 445 1 443  
2 446 1 443  
2 447 1 443  
2 448 1 443  
2 449 1 443  
2 450 1 443  
2 451 1 443  
2 452 1 443  
2 453 1 443  
2 454 1 443  
2 455 1 443  
2 456 1 443  
2 457 1 443  
2 458 1 443  
2 459 1 443  
1 460 0 16 0 
2 461 1 460  
2 462 1 460  
2 463 1 460  
2 464 1 460  
2 465 1 460  
2 466 1 460  
2 467 1 460  
2 468 1 460  
2 469 1 460  
2 470 1 460  
2 471 1 460  
2 472 1 460  
2 473 1 460  
2 474 1 460  
2 475 1 460  
2 476 1 460  
1 477 0 16 0 
2 478 1 477  
2 479 1 477  
2 480 1 477  
2 481 1 477  
2 482 1 477  
2 483 1 477  
2 484 1 477  
2 485 1 477  
2 486 1 477  
2 487 1 477  
2 488 1 477  
2 489 1 477  
2 490 1 477  
2 491 1 477  
2 492 1 477  
2 493 1 477  
1 494 0 16 0 
2 495 1 494  
2 496 1 494  
2 497 1 494  
2 498 1 494  
2 499 1 494  
2 500 1 494  
2 501 1 494  
2 502 1 494  
2 503 1 494  
2 504 1 494  
2 505 1 494  
2 506 1 494  
2 507 1 494  
2 508 1 494  
2 509 1 494  
2 510 1 494  
1 511 0 16 0 
2 512 1 511  
2 513 1 511  
2 514 1 511  
2 515 1 511  
2 516 1 511  
2 517 1 511  
2 518 1 511  
2 519 1 511  
2 520 1 511  
2 521 1 511  
2 522 1 511  
2 523 1 511  
2 524 1 511  
2 525 1 511  
2 526 1 511  
2 527 1 511  
1 528 0 16 0 
2 529 1 528  
2 530 1 528  
2 531 1 528  
2 532 1 528  
2 533 1 528  
2 534 1 528  
2 535 1 528  
2 536 1 528  
2 537 1 528  
2 538 1 528  
2 539 1 528  
2 540 1 528  
2 541 1 528  
2 542 1 528  
2 543 1 528  
2 544 1 528  
3 545 7 0 2 2 274 
0 546 7 2 2 3 291 
2 547 1 546  
2 548 1 546  
0 549 7 2 2 4 308 
2 550 1 549  
2 551 1 549  
0 552 7 2 2 5 325 
2 553 1 552  
2 554 1 552  
0 555 7 2 2 6 342 
2 556 1 555  
2 557 1 555  
0 558 7 2 2 7 359 
2 559 1 558  
2 560 1 558  
0 561 7 2 2 8 376 
2 562 1 561  
2 563 1 561  
0 564 7 2 2 9 393 
2 565 1 564  
2 566 1 564  
0 567 7 2 2 10 410 
2 568 1 567  
2 569 1 567  
0 570 7 2 2 11 427 
2 571 1 570  
2 572 1 570  
0 573 7 2 2 12 444 
2 574 1 573  
2 575 1 573  
0 576 7 2 2 13 461 
2 577 1 576  
2 578 1 576  
0 579 7 2 2 14 478 
2 580 1 579  
2 581 1 579  
0 582 7 2 2 15 495 
2 583 1 582  
2 584 1 582  
0 585 7 2 2 16 512 
2 586 1 585  
2 587 1 585  
0 588 7 2 2 17 529 
2 589 1 588  
2 590 1 588  
0 591 7 2 2 19 275 
2 592 1 591  
2 593 1 591  
0 594 7 2 2 20 292 
2 595 1 594  
2 596 1 594  
0 597 7 2 2 21 309 
2 598 1 597  
2 599 1 597  
0 600 7 2 2 22 326 
2 601 1 600  
2 602 1 600  
0 603 7 2 2 23 343 
2 604 1 603  
2 605 1 603  
0 606 7 2 2 24 360 
2 607 1 606  
2 608 1 606  
0 609 7 2 2 25 377 
2 610 1 609  
2 611 1 609  
0 612 7 2 2 26 394 
2 613 1 612  
2 614 1 612  
0 615 7 2 2 27 411 
2 616 1 615  
2 617 1 615  
0 618 7 2 2 28 428 
2 619 1 618  
2 620 1 618  
0 621 7 2 2 29 445 
2 622 1 621  
2 623 1 621  
0 624 7 2 2 30 462 
2 625 1 624  
2 626 1 624  
0 627 7 2 2 31 479 
2 628 1 627  
2 629 1 627  
0 630 7 2 2 32 496 
2 631 1 630  
2 632 1 630  
0 633 7 2 2 33 513 
2 634 1 633  
2 635 1 633  
0 636 7 2 2 34 530 
2 637 1 636  
2 638 1 636  
0 639 7 2 2 36 276 
2 640 1 639  
2 641 1 639  
0 642 7 2 2 37 293 
2 643 1 642  
2 644 1 642  
0 645 7 2 2 38 310 
2 646 1 645  
2 647 1 645  
0 648 7 2 2 39 327 
2 649 1 648  
2 650 1 648  
0 651 7 2 2 40 344 
2 652 1 651  
2 653 1 651  
0 654 7 2 2 41 361 
2 655 1 654  
2 656 1 654  
0 657 7 2 2 42 378 
2 658 1 657  
2 659 1 657  
0 660 7 2 2 43 395 
2 661 1 660  
2 662 1 660  
0 663 7 2 2 44 412 
2 664 1 663  
2 665 1 663  
0 666 7 2 2 45 429 
2 667 1 666  
2 668 1 666  
0 669 7 2 2 46 446 
2 670 1 669  
2 671 1 669  
0 672 7 2 2 47 463 
2 673 1 672  
2 674 1 672  
0 675 7 2 2 48 480 
2 676 1 675  
2 677 1 675  
0 678 7 2 2 49 497 
2 679 1 678  
2 680 1 678  
0 681 7 2 2 50 514 
2 682 1 681  
2 683 1 681  
0 684 7 2 2 51 531 
2 685 1 684  
2 686 1 684  
0 687 7 2 2 53 277 
2 688 1 687  
2 689 1 687  
0 690 7 2 2 54 294 
2 691 1 690  
2 692 1 690  
0 693 7 2 2 55 311 
2 694 1 693  
2 695 1 693  
0 696 7 2 2 56 328 
2 697 1 696  
2 698 1 696  
0 699 7 2 2 57 345 
2 700 1 699  
2 701 1 699  
0 702 7 2 2 58 362 
2 703 1 702  
2 704 1 702  
0 705 7 2 2 59 379 
2 706 1 705  
2 707 1 705  
0 708 7 2 2 60 396 
2 709 1 708  
2 710 1 708  
0 711 7 2 2 61 413 
2 712 1 711  
2 713 1 711  
0 714 7 2 2 62 430 
2 715 1 714  
2 716 1 714  
0 717 7 2 2 63 447 
2 718 1 717  
2 719 1 717  
0 720 7 2 2 64 464 
2 721 1 720  
2 722 1 720  
0 723 7 2 2 65 481 
2 724 1 723  
2 725 1 723  
0 726 7 2 2 66 498 
2 727 1 726  
2 728 1 726  
0 729 7 2 2 67 515 
2 730 1 729  
2 731 1 729  
0 732 7 2 2 68 532 
2 733 1 732  
2 734 1 732  
0 735 7 2 2 70 278 
2 736 1 735  
2 737 1 735  
0 738 7 2 2 71 295 
2 739 1 738  
2 740 1 738  
0 741 7 2 2 72 312 
2 742 1 741  
2 743 1 741  
0 744 7 2 2 73 329 
2 745 1 744  
2 746 1 744  
0 747 7 2 2 74 346 
2 748 1 747  
2 749 1 747  
0 750 7 2 2 75 363 
2 751 1 750  
2 752 1 750  
0 753 7 2 2 76 380 
2 754 1 753  
2 755 1 753  
0 756 7 2 2 77 397 
2 757 1 756  
2 758 1 756  
0 759 7 2 2 78 414 
2 760 1 759  
2 761 1 759  
0 762 7 2 2 79 431 
2 763 1 762  
2 764 1 762  
0 765 7 2 2 80 448 
2 766 1 765  
2 767 1 765  
0 768 7 2 2 81 465 
2 769 1 768  
2 770 1 768  
0 771 7 2 2 82 482 
2 772 1 771  
2 773 1 771  
0 774 7 2 2 83 499 
2 775 1 774  
2 776 1 774  
0 777 7 2 2 84 516 
2 778 1 777  
2 779 1 777  
0 780 7 2 2 85 533 
2 781 1 780  
2 782 1 780  
0 783 7 2 2 87 279 
2 784 1 783  
2 785 1 783  
0 786 7 2 2 88 296 
2 787 1 786  
2 788 1 786  
0 789 7 2 2 89 313 
2 790 1 789  
2 791 1 789  
0 792 7 2 2 90 330 
2 793 1 792  
2 794 1 792  
0 795 7 2 2 91 347 
2 796 1 795  
2 797 1 795  
0 798 7 2 2 92 364 
2 799 1 798  
2 800 1 798  
0 801 7 2 2 93 381 
2 802 1 801  
2 803 1 801  
0 804 7 2 2 94 398 
2 805 1 804  
2 806 1 804  
0 807 7 2 2 95 415 
2 808 1 807  
2 809 1 807  
0 810 7 2 2 96 432 
2 811 1 810  
2 812 1 810  
0 813 7 2 2 97 449 
2 814 1 813  
2 815 1 813  
0 816 7 2 2 98 466 
2 817 1 816  
2 818 1 816  
0 819 7 2 2 99 483 
2 820 1 819  
2 821 1 819  
0 822 7 2 2 100 500 
2 823 1 822  
2 824 1 822  
0 825 7 2 2 101 517 
2 826 1 825  
2 827 1 825  
0 828 7 2 2 102 534 
2 829 1 828  
2 830 1 828  
0 831 7 2 2 104 280 
2 832 1 831  
2 833 1 831  
0 834 7 2 2 105 297 
2 835 1 834  
2 836 1 834  
0 837 7 2 2 106 314 
2 838 1 837  
2 839 1 837  
0 840 7 2 2 107 331 
2 841 1 840  
2 842 1 840  
0 843 7 2 2 108 348 
2 844 1 843  
2 845 1 843  
0 846 7 2 2 109 365 
2 847 1 846  
2 848 1 846  
0 849 7 2 2 110 382 
2 850 1 849  
2 851 1 849  
0 852 7 2 2 111 399 
2 853 1 852  
2 854 1 852  
0 855 7 2 2 112 416 
2 856 1 855  
2 857 1 855  
0 858 7 2 2 113 433 
2 859 1 858  
2 860 1 858  
0 861 7 2 2 114 450 
2 862 1 861  
2 863 1 861  
0 864 7 2 2 115 467 
2 865 1 864  
2 866 1 864  
0 867 7 2 2 116 484 
2 868 1 867  
2 869 1 867  
0 870 7 2 2 117 501 
2 871 1 870  
2 872 1 870  
0 873 7 2 2 118 518 
2 874 1 873  
2 875 1 873  
0 876 7 2 2 119 535 
2 877 1 876  
2 878 1 876  
0 879 7 2 2 121 281 
2 880 1 879  
2 881 1 879  
0 882 7 2 2 122 298 
2 883 1 882  
2 884 1 882  
0 885 7 2 2 123 315 
2 886 1 885  
2 887 1 885  
0 888 7 2 2 124 332 
2 889 1 888  
2 890 1 888  
0 891 7 2 2 125 349 
2 892 1 891  
2 893 1 891  
0 894 7 2 2 126 366 
2 895 1 894  
2 896 1 894  
0 897 7 2 2 127 383 
2 898 1 897  
2 899 1 897  
0 900 7 2 2 128 400 
2 901 1 900  
2 902 1 900  
0 903 7 2 2 129 417 
2 904 1 903  
2 905 1 903  
0 906 7 2 2 130 434 
2 907 1 906  
2 908 1 906  
0 909 7 2 2 131 451 
2 910 1 909  
2 911 1 909  
0 912 7 2 2 132 468 
2 913 1 912  
2 914 1 912  
0 915 7 2 2 133 485 
2 916 1 915  
2 917 1 915  
0 918 7 2 2 134 502 
2 919 1 918  
2 920 1 918  
0 921 7 2 2 135 519 
2 922 1 921  
2 923 1 921  
0 924 7 2 2 136 536 
2 925 1 924  
2 926 1 924  
0 927 7 2 2 138 282 
2 928 1 927  
2 929 1 927  
0 930 7 2 2 139 299 
2 931 1 930  
2 932 1 930  
0 933 7 2 2 140 316 
2 934 1 933  
2 935 1 933  
0 936 7 2 2 141 333 
2 937 1 936  
2 938 1 936  
0 939 7 2 2 142 350 
2 940 1 939  
2 941 1 939  
0 942 7 2 2 143 367 
2 943 1 942  
2 944 1 942  
0 945 7 2 2 144 384 
2 946 1 945  
2 947 1 945  
0 948 7 2 2 145 401 
2 949 1 948  
2 950 1 948  
0 951 7 2 2 146 418 
2 952 1 951  
2 953 1 951  
0 954 7 2 2 147 435 
2 955 1 954  
2 956 1 954  
0 957 7 2 2 148 452 
2 958 1 957  
2 959 1 957  
0 960 7 2 2 149 469 
2 961 1 960  
2 962 1 960  
0 963 7 2 2 150 486 
2 964 1 963  
2 965 1 963  
0 966 7 2 2 151 503 
2 967 1 966  
2 968 1 966  
0 969 7 2 2 152 520 
2 970 1 969  
2 971 1 969  
0 972 7 2 2 153 537 
2 973 1 972  
2 974 1 972  
0 975 7 2 2 155 283 
2 976 1 975  
2 977 1 975  
0 978 7 2 2 156 300 
2 979 1 978  
2 980 1 978  
0 981 7 2 2 157 317 
2 982 1 981  
2 983 1 981  
0 984 7 2 2 158 334 
2 985 1 984  
2 986 1 984  
0 987 7 2 2 159 351 
2 988 1 987  
2 989 1 987  
0 990 7 2 2 160 368 
2 991 1 990  
2 992 1 990  
0 993 7 2 2 161 385 
2 994 1 993  
2 995 1 993  
0 996 7 2 2 162 402 
2 997 1 996  
2 998 1 996  
0 999 7 2 2 163 419 
2 1000 1 999  
2 1001 1 999  
0 1002 7 2 2 164 436 
2 1003 1 1002  
2 1004 1 1002  
0 1005 7 2 2 165 453 
2 1006 1 1005  
2 1007 1 1005  
0 1008 7 2 2 166 470 
2 1009 1 1008  
2 1010 1 1008  
0 1011 7 2 2 167 487 
2 1012 1 1011  
2 1013 1 1011  
0 1014 7 2 2 168 504 
2 1015 1 1014  
2 1016 1 1014  
0 1017 7 2 2 169 521 
2 1018 1 1017  
2 1019 1 1017  
0 1020 7 2 2 170 538 
2 1021 1 1020  
2 1022 1 1020  
0 1023 7 2 2 172 284 
2 1024 1 1023  
2 1025 1 1023  
0 1026 7 2 2 173 301 
2 1027 1 1026  
2 1028 1 1026  
0 1029 7 2 2 174 318 
2 1030 1 1029  
2 1031 1 1029  
0 1032 7 2 2 175 335 
2 1033 1 1032  
2 1034 1 1032  
0 1035 7 2 2 176 352 
2 1036 1 1035  
2 1037 1 1035  
0 1038 7 2 2 177 369 
2 1039 1 1038  
2 1040 1 1038  
0 1041 7 2 2 178 386 
2 1042 1 1041  
2 1043 1 1041  
0 1044 7 2 2 179 403 
2 1045 1 1044  
2 1046 1 1044  
0 1047 7 2 2 180 420 
2 1048 1 1047  
2 1049 1 1047  
0 1050 7 2 2 181 437 
2 1051 1 1050  
2 1052 1 1050  
0 1053 7 2 2 182 454 
2 1054 1 1053  
2 1055 1 1053  
0 1056 7 2 2 183 471 
2 1057 1 1056  
2 1058 1 1056  
0 1059 7 2 2 184 488 
2 1060 1 1059  
2 1061 1 1059  
0 1062 7 2 2 185 505 
2 1063 1 1062  
2 1064 1 1062  
0 1065 7 2 2 186 522 
2 1066 1 1065  
2 1067 1 1065  
0 1068 7 2 2 187 539 
2 1069 1 1068  
2 1070 1 1068  
0 1071 7 2 2 189 285 
2 1072 1 1071  
2 1073 1 1071  
0 1074 7 2 2 190 302 
2 1075 1 1074  
2 1076 1 1074  
0 1077 7 2 2 191 319 
2 1078 1 1077  
2 1079 1 1077  
0 1080 7 2 2 192 336 
2 1081 1 1080  
2 1082 1 1080  
0 1083 7 2 2 193 353 
2 1084 1 1083  
2 1085 1 1083  
0 1086 7 2 2 194 370 
2 1087 1 1086  
2 1088 1 1086  
0 1089 7 2 2 195 387 
2 1090 1 1089  
2 1091 1 1089  
0 1092 7 2 2 196 404 
2 1093 1 1092  
2 1094 1 1092  
0 1095 7 2 2 197 421 
2 1096 1 1095  
2 1097 1 1095  
0 1098 7 2 2 198 438 
2 1099 1 1098  
2 1100 1 1098  
0 1101 7 2 2 199 455 
2 1102 1 1101  
2 1103 1 1101  
0 1104 7 2 2 200 472 
2 1105 1 1104  
2 1106 1 1104  
0 1107 7 2 2 201 489 
2 1108 1 1107  
2 1109 1 1107  
0 1110 7 2 2 202 506 
2 1111 1 1110  
2 1112 1 1110  
0 1113 7 2 2 203 523 
2 1114 1 1113  
2 1115 1 1113  
0 1116 7 2 2 204 540 
2 1117 1 1116  
2 1118 1 1116  
0 1119 7 2 2 206 286 
2 1120 1 1119  
2 1121 1 1119  
0 1122 7 2 2 207 303 
2 1123 1 1122  
2 1124 1 1122  
0 1125 7 2 2 208 320 
2 1126 1 1125  
2 1127 1 1125  
0 1128 7 2 2 209 337 
2 1129 1 1128  
2 1130 1 1128  
0 1131 7 2 2 210 354 
2 1132 1 1131  
2 1133 1 1131  
0 1134 7 2 2 211 371 
2 1135 1 1134  
2 1136 1 1134  
0 1137 7 2 2 212 388 
2 1138 1 1137  
2 1139 1 1137  
0 1140 7 2 2 213 405 
2 1141 1 1140  
2 1142 1 1140  
0 1143 7 2 2 214 422 
2 1144 1 1143  
2 1145 1 1143  
0 1146 7 2 2 215 439 
2 1147 1 1146  
2 1148 1 1146  
0 1149 7 2 2 216 456 
2 1150 1 1149  
2 1151 1 1149  
0 1152 7 2 2 217 473 
2 1153 1 1152  
2 1154 1 1152  
0 1155 7 2 2 218 490 
2 1156 1 1155  
2 1157 1 1155  
0 1158 7 2 2 219 507 
2 1159 1 1158  
2 1160 1 1158  
0 1161 7 2 2 220 524 
2 1162 1 1161  
2 1163 1 1161  
0 1164 7 2 2 221 541 
2 1165 1 1164  
2 1166 1 1164  
0 1167 7 2 2 223 287 
2 1168 1 1167  
2 1169 1 1167  
0 1170 7 2 2 224 304 
2 1171 1 1170  
2 1172 1 1170  
0 1173 7 2 2 225 321 
2 1174 1 1173  
2 1175 1 1173  
0 1176 7 2 2 226 338 
2 1177 1 1176  
2 1178 1 1176  
0 1179 7 2 2 227 355 
2 1180 1 1179  
2 1181 1 1179  
0 1182 7 2 2 228 372 
2 1183 1 1182  
2 1184 1 1182  
0 1185 7 2 2 229 389 
2 1186 1 1185  
2 1187 1 1185  
0 1188 7 2 2 230 406 
2 1189 1 1188  
2 1190 1 1188  
0 1191 7 2 2 231 423 
2 1192 1 1191  
2 1193 1 1191  
0 1194 7 2 2 232 440 
2 1195 1 1194  
2 1196 1 1194  
0 1197 7 2 2 233 457 
2 1198 1 1197  
2 1199 1 1197  
0 1200 7 2 2 234 474 
2 1201 1 1200  
2 1202 1 1200  
0 1203 7 2 2 235 491 
2 1204 1 1203  
2 1205 1 1203  
0 1206 7 2 2 236 508 
2 1207 1 1206  
2 1208 1 1206  
0 1209 7 2 2 237 525 
2 1210 1 1209  
2 1211 1 1209  
0 1212 7 2 2 238 542 
2 1213 1 1212  
2 1214 1 1212  
0 1215 7 2 2 240 288 
2 1216 1 1215  
2 1217 1 1215  
0 1218 7 2 2 241 305 
2 1219 1 1218  
2 1220 1 1218  
0 1221 7 2 2 242 322 
2 1222 1 1221  
2 1223 1 1221  
0 1224 7 2 2 243 339 
2 1225 1 1224  
2 1226 1 1224  
0 1227 7 2 2 244 356 
2 1228 1 1227  
2 1229 1 1227  
0 1230 7 2 2 245 373 
2 1231 1 1230  
2 1232 1 1230  
0 1233 7 2 2 246 390 
2 1234 1 1233  
2 1235 1 1233  
0 1236 7 2 2 247 407 
2 1237 1 1236  
2 1238 1 1236  
0 1239 7 2 2 248 424 
2 1240 1 1239  
2 1241 1 1239  
0 1242 7 2 2 249 441 
2 1243 1 1242  
2 1244 1 1242  
0 1245 7 2 2 250 458 
2 1246 1 1245  
2 1247 1 1245  
0 1248 7 2 2 251 475 
2 1249 1 1248  
2 1250 1 1248  
0 1251 7 2 2 252 492 
2 1252 1 1251  
2 1253 1 1251  
0 1254 7 2 2 253 509 
2 1255 1 1254  
2 1256 1 1254  
0 1257 7 2 2 254 526 
2 1258 1 1257  
2 1259 1 1257  
0 1260 7 2 2 255 543 
2 1261 1 1260  
2 1262 1 1260  
0 1263 7 2 2 257 289 
2 1264 1 1263  
2 1265 1 1263  
0 1266 7 2 2 258 306 
2 1267 1 1266  
2 1268 1 1266  
0 1269 7 2 2 259 323 
2 1270 1 1269  
2 1271 1 1269  
0 1272 7 2 2 260 340 
2 1273 1 1272  
2 1274 1 1272  
0 1275 7 2 2 261 357 
2 1276 1 1275  
2 1277 1 1275  
0 1278 7 2 2 262 374 
2 1279 1 1278  
2 1280 1 1278  
0 1281 7 2 2 263 391 
2 1282 1 1281  
2 1283 1 1281  
0 1284 7 2 2 264 408 
2 1285 1 1284  
2 1286 1 1284  
0 1287 7 2 2 265 425 
2 1288 1 1287  
2 1289 1 1287  
0 1290 7 2 2 266 442 
2 1291 1 1290  
2 1292 1 1290  
0 1293 7 2 2 267 459 
2 1294 1 1293  
2 1295 1 1293  
0 1296 7 2 2 268 476 
2 1297 1 1296  
2 1298 1 1296  
0 1299 7 2 2 269 493 
2 1300 1 1299  
2 1301 1 1299  
0 1302 7 2 2 270 510 
2 1303 1 1302  
2 1304 1 1302  
0 1305 7 2 2 271 527 
2 1306 1 1305  
2 1307 1 1305  
0 1308 7 2 2 272 544 
2 1309 1 1308  
2 1310 1 1308  
0 1311 5 3 1 592 
2 1312 1 1311  
2 1313 1 1311  
2 1314 1 1311  
0 1315 5 3 1 640 
2 1316 1 1315  
2 1317 1 1315  
2 1318 1 1315  
0 1319 5 3 1 688 
2 1320 1 1319  
2 1321 1 1319  
2 1322 1 1319  
0 1323 5 3 1 736 
2 1324 1 1323  
2 1325 1 1323  
2 1326 1 1323  
0 1327 5 3 1 784 
2 1328 1 1327  
2 1329 1 1327  
2 1330 1 1327  
0 1331 5 3 1 832 
2 1332 1 1331  
2 1333 1 1331  
2 1334 1 1331  
0 1335 5 3 1 880 
2 1336 1 1335  
2 1337 1 1335  
2 1338 1 1335  
0 1339 5 3 1 928 
2 1340 1 1339  
2 1341 1 1339  
2 1342 1 1339  
0 1343 5 3 1 976 
2 1344 1 1343  
2 1345 1 1343  
2 1346 1 1343  
0 1347 5 3 1 1024 
2 1348 1 1347  
2 1349 1 1347  
2 1350 1 1347  
0 1351 5 3 1 1072 
2 1352 1 1351  
2 1353 1 1351  
2 1354 1 1351  
0 1355 5 3 1 1120 
2 1356 1 1355  
2 1357 1 1355  
2 1358 1 1355  
0 1359 5 3 1 1168 
2 1360 1 1359  
2 1361 1 1359  
2 1362 1 1359  
0 1363 5 3 1 1216 
2 1364 1 1363  
2 1365 1 1363  
2 1366 1 1363  
0 1367 5 3 1 1264 
2 1368 1 1367  
2 1369 1 1367  
2 1370 1 1367  
0 1371 4 1 2 593 1312 
0 1372 5 1 1 1313 
0 1373 4 1 2 641 1316 
0 1374 5 1 1 1317 
0 1375 4 1 2 689 1320 
0 1376 5 1 1 1321 
0 1377 4 1 2 737 1324 
0 1378 5 1 1 1325 
0 1379 4 1 2 785 1328 
0 1380 5 1 1 1329 
0 1381 4 1 2 833 1332 
0 1382 5 1 1 1333 
0 1383 4 1 2 881 1336 
0 1384 5 1 1 1337 
0 1385 4 1 2 929 1340 
0 1386 5 1 1 1341 
0 1387 4 1 2 977 1344 
0 1388 5 1 1 1345 
0 1389 4 1 2 1025 1348 
0 1390 5 1 1 1349 
0 1391 4 1 2 1073 1352 
0 1392 5 1 1 1353 
0 1393 4 1 2 1121 1356 
0 1394 5 1 1 1357 
0 1395 4 1 2 1169 1360 
0 1396 5 1 1 1361 
0 1397 4 1 2 1217 1364 
0 1398 5 1 1 1365 
0 1399 4 1 2 1265 1368 
0 1400 5 1 1 1369 
0 1401 4 2 2 1371 1372 
2 1402 1 1401  
2 1403 1 1401  
0 1404 4 2 2 1373 1374 
2 1405 1 1404  
2 1406 1 1404  
0 1407 4 2 2 1375 1376 
2 1408 1 1407  
2 1409 1 1407  
0 1410 4 2 2 1377 1378 
2 1411 1 1410  
2 1412 1 1410  
0 1413 4 2 2 1379 1380 
2 1414 1 1413  
2 1415 1 1413  
0 1416 4 2 2 1381 1382 
2 1417 1 1416  
2 1418 1 1416  
0 1419 4 2 2 1383 1384 
2 1420 1 1419  
2 1421 1 1419  
0 1422 4 2 2 1385 1386 
2 1423 1 1422  
2 1424 1 1422  
0 1425 4 2 2 1387 1388 
2 1426 1 1425  
2 1427 1 1425  
0 1428 4 2 2 1389 1390 
2 1429 1 1428  
2 1430 1 1428  
0 1431 4 2 2 1391 1392 
2 1432 1 1431  
2 1433 1 1431  
0 1434 4 2 2 1393 1394 
2 1435 1 1434  
2 1436 1 1434  
0 1437 4 2 2 1395 1396 
2 1438 1 1437  
2 1439 1 1437  
0 1440 4 2 2 1397 1398 
2 1441 1 1440  
2 1442 1 1440  
0 1443 4 2 2 1399 1400 
2 1444 1 1443  
2 1445 1 1443  
0 1446 4 3 2 1402 547 
2 1447 1 1446  
2 1448 1 1446  
2 1449 1 1446  
0 1450 4 3 2 1405 595 
2 1451 1 1450  
2 1452 1 1450  
2 1453 1 1450  
0 1454 4 3 2 1408 643 
2 1455 1 1454  
2 1456 1 1454  
2 1457 1 1454  
0 1458 4 3 2 1411 691 
2 1459 1 1458  
2 1460 1 1458  
2 1461 1 1458  
0 1462 4 3 2 1414 739 
2 1463 1 1462  
2 1464 1 1462  
2 1465 1 1462  
0 1466 4 3 2 1417 787 
2 1467 1 1466  
2 1468 1 1466  
2 1469 1 1466  
0 1470 4 3 2 1420 835 
2 1471 1 1470  
2 1472 1 1470  
2 1473 1 1470  
0 1474 4 3 2 1423 883 
2 1475 1 1474  
2 1476 1 1474  
2 1477 1 1474  
0 1478 4 3 2 1426 931 
2 1479 1 1478  
2 1480 1 1478  
2 1481 1 1478  
0 1482 4 3 2 1429 979 
2 1483 1 1482  
2 1484 1 1482  
2 1485 1 1482  
0 1486 4 3 2 1432 1027 
2 1487 1 1486  
2 1488 1 1486  
2 1489 1 1486  
0 1490 4 3 2 1435 1075 
2 1491 1 1490  
2 1492 1 1490  
2 1493 1 1490  
0 1494 4 3 2 1438 1123 
2 1495 1 1494  
2 1496 1 1494  
2 1497 1 1494  
0 1498 4 3 2 1441 1171 
2 1499 1 1498  
2 1500 1 1498  
2 1501 1 1498  
0 1502 4 3 2 1444 1219 
2 1503 1 1502  
2 1504 1 1502  
2 1505 1 1502  
0 1506 4 1 2 1403 1447 
0 1507 4 1 2 1448 548 
0 1508 4 2 2 1314 1449 
2 1509 1 1508  
2 1510 1 1508  
0 1511 4 1 2 1406 1451 
0 1512 4 1 2 1452 596 
0 1513 4 2 2 1318 1453 
2 1514 1 1513  
2 1515 1 1513  
0 1516 4 1 2 1409 1455 
0 1517 4 1 2 1456 644 
0 1518 4 2 2 1322 1457 
2 1519 1 1518  
2 1520 1 1518  
0 1521 4 1 2 1412 1459 
0 1522 4 1 2 1460 692 
0 1523 4 2 2 1326 1461 
2 1524 1 1523  
2 1525 1 1523  
0 1526 4 1 2 1415 1463 
0 1527 4 1 2 1464 740 
0 1528 4 2 2 1330 1465 
2 1529 1 1528  
2 1530 1 1528  
0 1531 4 1 2 1418 1467 
0 1532 4 1 2 1468 788 
0 1533 4 2 2 1334 1469 
2 1534 1 1533  
2 1535 1 1533  
0 1536 4 1 2 1421 1471 
0 1537 4 1 2 1472 836 
0 1538 4 2 2 1338 1473 
2 1539 1 1538  
2 1540 1 1538  
0 1541 4 1 2 1424 1475 
0 1542 4 1 2 1476 884 
0 1543 4 2 2 1342 1477 
2 1544 1 1543  
2 1545 1 1543  
0 1546 4 1 2 1427 1479 
0 1547 4 1 2 1480 932 
0 1548 4 2 2 1346 1481 
2 1549 1 1548  
2 1550 1 1548  
0 1551 4 1 2 1430 1483 
0 1552 4 1 2 1484 980 
0 1553 4 2 2 1350 1485 
2 1554 1 1553  
2 1555 1 1553  
0 1556 4 1 2 1433 1487 
0 1557 4 1 2 1488 1028 
0 1558 4 2 2 1354 1489 
2 1559 1 1558  
2 1560 1 1558  
0 1561 4 1 2 1436 1491 
0 1562 4 1 2 1492 1076 
0 1563 4 2 2 1358 1493 
2 1564 1 1563  
2 1565 1 1563  
0 1566 4 1 2 1439 1495 
0 1567 4 1 2 1496 1124 
0 1568 4 2 2 1362 1497 
2 1569 1 1568  
2 1570 1 1568  
0 1571 4 1 2 1442 1499 
0 1572 4 1 2 1500 1172 
0 1573 4 2 2 1366 1501 
2 1574 1 1573  
2 1575 1 1573  
0 1576 4 1 2 1445 1503 
0 1577 4 1 2 1504 1220 
0 1578 4 2 2 1370 1505 
2 1579 1 1578  
2 1580 1 1578  
3 1581 4 0 2 1506 1507 
0 1582 4 2 2 1511 1512 
2 1583 1 1582  
2 1584 1 1582  
0 1585 4 2 2 1516 1517 
2 1586 1 1585  
2 1587 1 1585  
0 1588 4 2 2 1521 1522 
2 1589 1 1588  
2 1590 1 1588  
0 1591 4 2 2 1526 1527 
2 1592 1 1591  
2 1593 1 1591  
0 1594 4 2 2 1531 1532 
2 1595 1 1594  
2 1596 1 1594  
0 1597 4 2 2 1536 1537 
2 1598 1 1597  
2 1599 1 1597  
0 1600 4 2 2 1541 1542 
2 1601 1 1600  
2 1602 1 1600  
0 1603 4 2 2 1546 1547 
2 1604 1 1603  
2 1605 1 1603  
0 1606 4 2 2 1551 1552 
2 1607 1 1606  
2 1608 1 1606  
0 1609 4 2 2 1556 1557 
2 1610 1 1609  
2 1611 1 1609  
0 1612 4 2 2 1561 1562 
2 1613 1 1612  
2 1614 1 1612  
0 1615 4 2 2 1566 1567 
2 1616 1 1615  
2 1617 1 1615  
0 1618 4 2 2 1571 1572 
2 1619 1 1618  
2 1620 1 1618  
0 1621 4 2 2 1576 1577 
2 1622 1 1621  
2 1623 1 1621  
0 1624 4 3 2 1267 1579 
2 1625 1 1624  
2 1626 1 1624  
2 1627 1 1624  
0 1628 4 3 2 1583 1509 
2 1629 1 1628  
2 1630 1 1628  
2 1631 1 1628  
0 1632 4 3 2 1586 1514 
2 1633 1 1632  
2 1634 1 1632  
2 1635 1 1632  
0 1636 4 3 2 1589 1519 
2 1637 1 1636  
2 1638 1 1636  
2 1639 1 1636  
0 1640 4 3 2 1592 1524 
2 1641 1 1640  
2 1642 1 1640  
2 1643 1 1640  
0 1644 4 3 2 1595 1529 
2 1645 1 1644  
2 1646 1 1644  
2 1647 1 1644  
0 1648 4 3 2 1598 1534 
2 1649 1 1648  
2 1650 1 1648  
2 1651 1 1648  
0 1652 4 3 2 1601 1539 
2 1653 1 1652  
2 1654 1 1652  
2 1655 1 1652  
0 1656 4 3 2 1604 1544 
2 1657 1 1656  
2 1658 1 1656  
2 1659 1 1656  
0 1660 4 3 2 1607 1549 
2 1661 1 1660  
2 1662 1 1660  
2 1663 1 1660  
0 1664 4 3 2 1610 1554 
2 1665 1 1664  
2 1666 1 1664  
2 1667 1 1664  
0 1668 4 3 2 1613 1559 
2 1669 1 1668  
2 1670 1 1668  
2 1671 1 1668  
0 1672 4 3 2 1616 1564 
2 1673 1 1672  
2 1674 1 1672  
2 1675 1 1672  
0 1676 4 3 2 1619 1569 
2 1677 1 1676  
2 1678 1 1676  
2 1679 1 1676  
0 1680 4 3 2 1622 1574 
2 1681 1 1680  
2 1682 1 1680  
2 1683 1 1680  
0 1684 4 1 2 1268 1625 
0 1685 4 1 2 1626 1580 
0 1686 4 1 2 1584 1629 
0 1687 4 1 2 1630 1510 
0 1688 4 1 2 1587 1633 
0 1689 4 1 2 1634 1515 
0 1690 4 1 2 1590 1637 
0 1691 4 1 2 1638 1520 
0 1692 4 1 2 1593 1641 
0 1693 4 1 2 1642 1525 
0 1694 4 1 2 1596 1645 
0 1695 4 1 2 1646 1530 
0 1696 4 1 2 1599 1649 
0 1697 4 1 2 1650 1535 
0 1698 4 1 2 1602 1653 
0 1699 4 1 2 1654 1540 
0 1700 4 1 2 1605 1657 
0 1701 4 1 2 1658 1545 
0 1702 4 1 2 1608 1661 
0 1703 4 1 2 1662 1550 
0 1704 4 1 2 1611 1665 
0 1705 4 1 2 1666 1555 
0 1706 4 1 2 1614 1669 
0 1707 4 1 2 1670 1560 
0 1708 4 1 2 1617 1673 
0 1709 4 1 2 1674 1565 
0 1710 4 1 2 1620 1677 
0 1711 4 1 2 1678 1570 
0 1712 4 1 2 1623 1681 
0 1713 4 1 2 1682 1575 
0 1714 4 2 2 1684 1685 
2 1715 1 1714  
2 1716 1 1714  
0 1717 4 2 2 1686 1687 
2 1718 1 1717  
2 1719 1 1717  
0 1720 4 2 2 1688 1689 
2 1721 1 1720  
2 1722 1 1720  
0 1723 4 2 2 1690 1691 
2 1724 1 1723  
2 1725 1 1723  
0 1726 4 2 2 1692 1693 
2 1727 1 1726  
2 1728 1 1726  
0 1729 4 2 2 1694 1695 
2 1730 1 1729  
2 1731 1 1729  
0 1732 4 2 2 1696 1697 
2 1733 1 1732  
2 1734 1 1732  
0 1735 4 2 2 1698 1699 
2 1736 1 1735  
2 1737 1 1735  
0 1738 4 2 2 1700 1701 
2 1739 1 1738  
2 1740 1 1738  
0 1741 4 2 2 1702 1703 
2 1742 1 1741  
2 1743 1 1741  
0 1744 4 2 2 1704 1705 
2 1745 1 1744  
2 1746 1 1744  
0 1747 4 2 2 1706 1707 
2 1748 1 1747  
2 1749 1 1747  
0 1750 4 2 2 1708 1709 
2 1751 1 1750  
2 1752 1 1750  
0 1753 4 2 2 1710 1711 
2 1754 1 1753  
2 1755 1 1753  
0 1756 4 2 2 1712 1713 
2 1757 1 1756  
2 1758 1 1756  
0 1759 4 3 2 1715 1222 
2 1760 1 1759  
2 1761 1 1759  
2 1762 1 1759  
0 1763 4 3 2 1718 550 
2 1764 1 1763  
2 1765 1 1763  
2 1766 1 1763  
0 1767 4 3 2 1721 598 
2 1768 1 1767  
2 1769 1 1767  
2 1770 1 1767  
0 1771 4 3 2 1724 646 
2 1772 1 1771  
2 1773 1 1771  
2 1774 1 1771  
0 1775 4 3 2 1727 694 
2 1776 1 1775  
2 1777 1 1775  
2 1778 1 1775  
0 1779 4 3 2 1730 742 
2 1780 1 1779  
2 1781 1 1779  
2 1782 1 1779  
0 1783 4 3 2 1733 790 
2 1784 1 1783  
2 1785 1 1783  
2 1786 1 1783  
0 1787 4 3 2 1736 838 
2 1788 1 1787  
2 1789 1 1787  
2 1790 1 1787  
0 1791 4 3 2 1739 886 
2 1792 1 1791  
2 1793 1 1791  
2 1794 1 1791  
0 1795 4 3 2 1742 934 
2 1796 1 1795  
2 1797 1 1795  
2 1798 1 1795  
0 1799 4 3 2 1745 982 
2 1800 1 1799  
2 1801 1 1799  
2 1802 1 1799  
0 1803 4 3 2 1748 1030 
2 1804 1 1803  
2 1805 1 1803  
2 1806 1 1803  
0 1807 4 3 2 1751 1078 
2 1808 1 1807  
2 1809 1 1807  
2 1810 1 1807  
0 1811 4 3 2 1754 1126 
2 1812 1 1811  
2 1813 1 1811  
2 1814 1 1811  
0 1815 4 3 2 1757 1174 
2 1816 1 1815  
2 1817 1 1815  
2 1818 1 1815  
0 1819 4 1 2 1716 1760 
0 1820 4 1 2 1761 1223 
0 1821 4 2 2 1627 1762 
2 1822 1 1821  
2 1823 1 1821  
0 1824 4 1 2 1719 1764 
0 1825 4 1 2 1765 551 
0 1826 4 2 2 1631 1766 
2 1827 1 1826  
2 1828 1 1826  
0 1829 4 1 2 1722 1768 
0 1830 4 1 2 1769 599 
0 1831 4 2 2 1635 1770 
2 1832 1 1831  
2 1833 1 1831  
0 1834 4 1 2 1725 1772 
0 1835 4 1 2 1773 647 
0 1836 4 2 2 1639 1774 
2 1837 1 1836  
2 1838 1 1836  
0 1839 4 1 2 1728 1776 
0 1840 4 1 2 1777 695 
0 1841 4 2 2 1643 1778 
2 1842 1 1841  
2 1843 1 1841  
0 1844 4 1 2 1731 1780 
0 1845 4 1 2 1781 743 
0 1846 4 2 2 1647 1782 
2 1847 1 1846  
2 1848 1 1846  
0 1849 4 1 2 1734 1784 
0 1850 4 1 2 1785 791 
0 1851 4 2 2 1651 1786 
2 1852 1 1851  
2 1853 1 1851  
0 1854 4 1 2 1737 1788 
0 1855 4 1 2 1789 839 
0 1856 4 2 2 1655 1790 
2 1857 1 1856  
2 1858 1 1856  
0 1859 4 1 2 1740 1792 
0 1860 4 1 2 1793 887 
0 1861 4 2 2 1659 1794 
2 1862 1 1861  
2 1863 1 1861  
0 1864 4 1 2 1743 1796 
0 1865 4 1 2 1797 935 
0 1866 4 2 2 1663 1798 
2 1867 1 1866  
2 1868 1 1866  
0 1869 4 1 2 1746 1800 
0 1870 4 1 2 1801 983 
0 1871 4 2 2 1667 1802 
2 1872 1 1871  
2 1873 1 1871  
0 1874 4 1 2 1749 1804 
0 1875 4 1 2 1805 1031 
0 1876 4 2 2 1671 1806 
2 1877 1 1876  
2 1878 1 1876  
0 1879 4 1 2 1752 1808 
0 1880 4 1 2 1809 1079 
0 1881 4 2 2 1675 1810 
2 1882 1 1881  
2 1883 1 1881  
0 1884 4 1 2 1755 1812 
0 1885 4 1 2 1813 1127 
0 1886 4 2 2 1679 1814 
2 1887 1 1886  
2 1888 1 1886  
0 1889 4 1 2 1758 1816 
0 1890 4 1 2 1817 1175 
0 1891 4 2 2 1683 1818 
2 1892 1 1891  
2 1893 1 1891  
0 1894 4 2 2 1819 1820 
2 1895 1 1894  
2 1896 1 1894  
0 1897 4 3 2 1270 1822 
2 1898 1 1897  
2 1899 1 1897  
2 1900 1 1897  
3 1901 4 0 2 1824 1825 
0 1902 4 2 2 1829 1830 
2 1903 1 1902  
2 1904 1 1902  
0 1905 4 2 2 1834 1835 
2 1906 1 1905  
2 1907 1 1905  
0 1908 4 2 2 1839 1840 
2 1909 1 1908  
2 1910 1 1908  
0 1911 4 2 2 1844 1845 
2 1912 1 1911  
2 1913 1 1911  
0 1914 4 2 2 1849 1850 
2 1915 1 1914  
2 1916 1 1914  
0 1917 4 2 2 1854 1855 
2 1918 1 1917  
2 1919 1 1917  
0 1920 4 2 2 1859 1860 
2 1921 1 1920  
2 1922 1 1920  
0 1923 4 2 2 1864 1865 
2 1924 1 1923  
2 1925 1 1923  
0 1926 4 2 2 1869 1870 
2 1927 1 1926  
2 1928 1 1926  
0 1929 4 2 2 1874 1875 
2 1930 1 1929  
2 1931 1 1929  
0 1932 4 2 2 1879 1880 
2 1933 1 1932  
2 1934 1 1932  
0 1935 4 2 2 1884 1885 
2 1936 1 1935  
2 1937 1 1935  
0 1938 4 2 2 1889 1890 
2 1939 1 1938  
2 1940 1 1938  
0 1941 4 3 2 1895 1892 
2 1942 1 1941  
2 1943 1 1941  
2 1944 1 1941  
0 1945 4 1 2 1271 1898 
0 1946 4 1 2 1899 1823 
0 1947 4 3 2 1903 1827 
2 1948 1 1947  
2 1949 1 1947  
2 1950 1 1947  
0 1951 4 3 2 1906 1832 
2 1952 1 1951  
2 1953 1 1951  
2 1954 1 1951  
0 1955 4 3 2 1909 1837 
2 1956 1 1955  
2 1957 1 1955  
2 1958 1 1955  
0 1959 4 3 2 1912 1842 
2 1960 1 1959  
2 1961 1 1959  
2 1962 1 1959  
0 1963 4 3 2 1915 1847 
2 1964 1 1963  
2 1965 1 1963  
2 1966 1 1963  
0 1967 4 3 2 1918 1852 
2 1968 1 1967  
2 1969 1 1967  
2 1970 1 1967  
0 1971 4 3 2 1921 1857 
2 1972 1 1971  
2 1973 1 1971  
2 1974 1 1971  
0 1975 4 3 2 1924 1862 
2 1976 1 1975  
2 1977 1 1975  
2 1978 1 1975  
0 1979 4 3 2 1927 1867 
2 1980 1 1979  
2 1981 1 1979  
2 1982 1 1979  
0 1983 4 3 2 1930 1872 
2 1984 1 1983  
2 1985 1 1983  
2 1986 1 1983  
0 1987 4 3 2 1933 1877 
2 1988 1 1987  
2 1989 1 1987  
2 1990 1 1987  
0 1991 4 3 2 1936 1882 
2 1992 1 1991  
2 1993 1 1991  
2 1994 1 1991  
0 1995 4 3 2 1939 1887 
2 1996 1 1995  
2 1997 1 1995  
2 1998 1 1995  
0 1999 4 1 2 1896 1942 
0 2000 4 1 2 1943 1893 
0 2001 4 2 2 1945 1946 
2 2002 1 2001  
2 2003 1 2001  
0 2004 4 1 2 1904 1948 
0 2005 4 1 2 1949 1828 
0 2006 4 1 2 1907 1952 
0 2007 4 1 2 1953 1833 
0 2008 4 1 2 1910 1956 
0 2009 4 1 2 1957 1838 
0 2010 4 1 2 1913 1960 
0 2011 4 1 2 1961 1843 
0 2012 4 1 2 1916 1964 
0 2013 4 1 2 1965 1848 
0 2014 4 1 2 1919 1968 
0 2015 4 1 2 1969 1853 
0 2016 4 1 2 1922 1972 
0 2017 4 1 2 1973 1858 
0 2018 4 1 2 1925 1976 
0 2019 4 1 2 1977 1863 
0 2020 4 1 2 1928 1980 
0 2021 4 1 2 1981 1868 
0 2022 4 1 2 1931 1984 
0 2023 4 1 2 1985 1873 
0 2024 4 1 2 1934 1988 
0 2025 4 1 2 1989 1878 
0 2026 4 1 2 1937 1992 
0 2027 4 1 2 1993 1883 
0 2028 4 1 2 1940 1996 
0 2029 4 1 2 1997 1888 
0 2030 4 2 2 1999 2000 
2 2031 1 2030  
2 2032 1 2030  
0 2033 4 3 2 2002 1225 
2 2034 1 2033  
2 2035 1 2033  
2 2036 1 2033  
0 2037 4 2 2 2004 2005 
2 2038 1 2037  
2 2039 1 2037  
0 2040 4 2 2 2006 2007 
2 2041 1 2040  
2 2042 1 2040  
0 2043 4 2 2 2008 2009 
2 2044 1 2043  
2 2045 1 2043  
0 2046 4 2 2 2010 2011 
2 2047 1 2046  
2 2048 1 2046  
0 2049 4 2 2 2012 2013 
2 2050 1 2049  
2 2051 1 2049  
0 2052 4 2 2 2014 2015 
2 2053 1 2052  
2 2054 1 2052  
0 2055 4 2 2 2016 2017 
2 2056 1 2055  
2 2057 1 2055  
0 2058 4 2 2 2018 2019 
2 2059 1 2058  
2 2060 1 2058  
0 2061 4 2 2 2020 2021 
2 2062 1 2061  
2 2063 1 2061  
0 2064 4 2 2 2022 2023 
2 2065 1 2064  
2 2066 1 2064  
0 2067 4 2 2 2024 2025 
2 2068 1 2067  
2 2069 1 2067  
0 2070 4 2 2 2026 2027 
2 2071 1 2070  
2 2072 1 2070  
0 2073 4 2 2 2028 2029 
2 2074 1 2073  
2 2075 1 2073  
0 2076 4 3 2 2031 1177 
2 2077 1 2076  
2 2078 1 2076  
2 2079 1 2076  
0 2080 4 1 2 2003 2034 
0 2081 4 1 2 2035 1226 
0 2082 4 2 2 1900 2036 
2 2083 1 2082  
2 2084 1 2082  
0 2085 4 3 2 2038 553 
2 2086 1 2085  
2 2087 1 2085  
2 2088 1 2085  
0 2089 4 3 2 2041 601 
2 2090 1 2089  
2 2091 1 2089  
2 2092 1 2089  
0 2093 4 3 2 2044 649 
2 2094 1 2093  
2 2095 1 2093  
2 2096 1 2093  
0 2097 4 3 2 2047 697 
2 2098 1 2097  
2 2099 1 2097  
2 2100 1 2097  
0 2101 4 3 2 2050 745 
2 2102 1 2101  
2 2103 1 2101  
2 2104 1 2101  
0 2105 4 3 2 2053 793 
2 2106 1 2105  
2 2107 1 2105  
2 2108 1 2105  
0 2109 4 3 2 2056 841 
2 2110 1 2109  
2 2111 1 2109  
2 2112 1 2109  
0 2113 4 3 2 2059 889 
2 2114 1 2113  
2 2115 1 2113  
2 2116 1 2113  
0 2117 4 3 2 2062 937 
2 2118 1 2117  
2 2119 1 2117  
2 2120 1 2117  
0 2121 4 3 2 2065 985 
2 2122 1 2121  
2 2123 1 2121  
2 2124 1 2121  
0 2125 4 3 2 2068 1033 
2 2126 1 2125  
2 2127 1 2125  
2 2128 1 2125  
0 2129 4 3 2 2071 1081 
2 2130 1 2129  
2 2131 1 2129  
2 2132 1 2129  
0 2133 4 3 2 2074 1129 
2 2134 1 2133  
2 2135 1 2133  
2 2136 1 2133  
0 2137 4 1 2 2032 2077 
0 2138 4 1 2 2078 1178 
0 2139 4 2 2 1944 2079 
2 2140 1 2139  
2 2141 1 2139  
0 2142 4 2 2 2080 2081 
2 2143 1 2142  
2 2144 1 2142  
0 2145 4 3 2 1273 2083 
2 2146 1 2145  
2 2147 1 2145  
2 2148 1 2145  
0 2149 4 1 2 2039 2086 
0 2150 4 1 2 2087 554 
0 2151 4 2 2 1950 2088 
2 2152 1 2151  
2 2153 1 2151  
0 2154 4 1 2 2042 2090 
0 2155 4 1 2 2091 602 
0 2156 4 2 2 1954 2092 
2 2157 1 2156  
2 2158 1 2156  
0 2159 4 1 2 2045 2094 
0 2160 4 1 2 2095 650 
0 2161 4 2 2 1958 2096 
2 2162 1 2161  
2 2163 1 2161  
0 2164 4 1 2 2048 2098 
0 2165 4 1 2 2099 698 
0 2166 4 2 2 1962 2100 
2 2167 1 2166  
2 2168 1 2166  
0 2169 4 1 2 2051 2102 
0 2170 4 1 2 2103 746 
0 2171 4 2 2 1966 2104 
2 2172 1 2171  
2 2173 1 2171  
0 2174 4 1 2 2054 2106 
0 2175 4 1 2 2107 794 
0 2176 4 2 2 1970 2108 
2 2177 1 2176  
2 2178 1 2176  
0 2179 4 1 2 2057 2110 
0 2180 4 1 2 2111 842 
0 2181 4 2 2 1974 2112 
2 2182 1 2181  
2 2183 1 2181  
0 2184 4 1 2 2060 2114 
0 2185 4 1 2 2115 890 
0 2186 4 2 2 1978 2116 
2 2187 1 2186  
2 2188 1 2186  
0 2189 4 1 2 2063 2118 
0 2190 4 1 2 2119 938 
0 2191 4 2 2 1982 2120 
2 2192 1 2191  
2 2193 1 2191  
0 2194 4 1 2 2066 2122 
0 2195 4 1 2 2123 986 
0 2196 4 2 2 1986 2124 
2 2197 1 2196  
2 2198 1 2196  
0 2199 4 1 2 2069 2126 
0 2200 4 1 2 2127 1034 
0 2201 4 2 2 1990 2128 
2 2202 1 2201  
2 2203 1 2201  
0 2204 4 1 2 2072 2130 
0 2205 4 1 2 2131 1082 
0 2206 4 2 2 1994 2132 
2 2207 1 2206  
2 2208 1 2206  
0 2209 4 1 2 2075 2134 
0 2210 4 1 2 2135 1130 
0 2211 4 2 2 1998 2136 
2 2212 1 2211  
2 2213 1 2211  
0 2214 4 2 2 2137 2138 
2 2215 1 2214  
2 2216 1 2214  
0 2217 4 3 2 2143 2140 
2 2218 1 2217  
2 2219 1 2217  
2 2220 1 2217  
0 2221 4 1 2 1274 2146 
0 2222 4 1 2 2147 2084 
3 2223 4 0 2 2149 2150 
0 2224 4 2 2 2154 2155 
2 2225 1 2224  
2 2226 1 2224  
0 2227 4 2 2 2159 2160 
2 2228 1 2227  
2 2229 1 2227  
0 2230 4 2 2 2164 2165 
2 2231 1 2230  
2 2232 1 2230  
0 2233 4 2 2 2169 2170 
2 2234 1 2233  
2 2235 1 2233  
0 2236 4 2 2 2174 2175 
2 2237 1 2236  
2 2238 1 2236  
0 2239 4 2 2 2179 2180 
2 2240 1 2239  
2 2241 1 2239  
0 2242 4 2 2 2184 2185 
2 2243 1 2242  
2 2244 1 2242  
0 2245 4 2 2 2189 2190 
2 2246 1 2245  
2 2247 1 2245  
0 2248 4 2 2 2194 2195 
2 2249 1 2248  
2 2250 1 2248  
0 2251 4 2 2 2199 2200 
2 2252 1 2251  
2 2253 1 2251  
0 2254 4 2 2 2204 2205 
2 2255 1 2254  
2 2256 1 2254  
0 2257 4 2 2 2209 2210 
2 2258 1 2257  
2 2259 1 2257  
0 2260 4 3 2 2215 2212 
2 2261 1 2260  
2 2262 1 2260  
2 2263 1 2260  
0 2264 4 1 2 2144 2218 
0 2265 4 1 2 2219 2141 
0 2266 4 2 2 2221 2222 
2 2267 1 2266  
2 2268 1 2266  
0 2269 4 3 2 2225 2152 
2 2270 1 2269  
2 2271 1 2269  
2 2272 1 2269  
0 2273 4 3 2 2228 2157 
2 2274 1 2273  
2 2275 1 2273  
2 2276 1 2273  
0 2277 4 3 2 2231 2162 
2 2278 1 2277  
2 2279 1 2277  
2 2280 1 2277  
0 2281 4 3 2 2234 2167 
2 2282 1 2281  
2 2283 1 2281  
2 2284 1 2281  
0 2285 4 3 2 2237 2172 
2 2286 1 2285  
2 2287 1 2285  
2 2288 1 2285  
0 2289 4 3 2 2240 2177 
2 2290 1 2289  
2 2291 1 2289  
2 2292 1 2289  
0 2293 4 3 2 2243 2182 
2 2294 1 2293  
2 2295 1 2293  
2 2296 1 2293  
0 2297 4 3 2 2246 2187 
2 2298 1 2297  
2 2299 1 2297  
2 2300 1 2297  
0 2301 4 3 2 2249 2192 
2 2302 1 2301  
2 2303 1 2301  
2 2304 1 2301  
0 2305 4 3 2 2252 2197 
2 2306 1 2305  
2 2307 1 2305  
2 2308 1 2305  
0 2309 4 3 2 2255 2202 
2 2310 1 2309  
2 2311 1 2309  
2 2312 1 2309  
0 2313 4 3 2 2258 2207 
2 2314 1 2313  
2 2315 1 2313  
2 2316 1 2313  
0 2317 4 1 2 2216 2261 
0 2318 4 1 2 2262 2213 
0 2319 4 2 2 2264 2265 
2 2320 1 2319  
2 2321 1 2319  
0 2322 4 3 2 2267 1228 
2 2323 1 2322  
2 2324 1 2322  
2 2325 1 2322  
0 2326 4 1 2 2226 2270 
0 2327 4 1 2 2271 2153 
0 2328 4 1 2 2229 2274 
0 2329 4 1 2 2275 2158 
0 2330 4 1 2 2232 2278 
0 2331 4 1 2 2279 2163 
0 2332 4 1 2 2235 2282 
0 2333 4 1 2 2283 2168 
0 2334 4 1 2 2238 2286 
0 2335 4 1 2 2287 2173 
0 2336 4 1 2 2241 2290 
0 2337 4 1 2 2291 2178 
0 2338 4 1 2 2244 2294 
0 2339 4 1 2 2295 2183 
0 2340 4 1 2 2247 2298 
0 2341 4 1 2 2299 2188 
0 2342 4 1 2 2250 2302 
0 2343 4 1 2 2303 2193 
0 2344 4 1 2 2253 2306 
0 2345 4 1 2 2307 2198 
0 2346 4 1 2 2256 2310 
0 2347 4 1 2 2311 2203 
0 2348 4 1 2 2259 2314 
0 2349 4 1 2 2315 2208 
0 2350 4 2 2 2317 2318 
2 2351 1 2350  
2 2352 1 2350  
0 2353 4 3 2 2320 1180 
2 2354 1 2353  
2 2355 1 2353  
2 2356 1 2353  
0 2357 4 1 2 2268 2323 
0 2358 4 1 2 2324 1229 
0 2359 4 2 2 2148 2325 
2 2360 1 2359  
2 2361 1 2359  
0 2362 4 2 2 2326 2327 
2 2363 1 2362  
2 2364 1 2362  
0 2365 4 2 2 2328 2329 
2 2366 1 2365  
2 2367 1 2365  
0 2368 4 2 2 2330 2331 
2 2369 1 2368  
2 2370 1 2368  
0 2371 4 2 2 2332 2333 
2 2372 1 2371  
2 2373 1 2371  
0 2374 4 2 2 2334 2335 
2 2375 1 2374  
2 2376 1 2374  
0 2377 4 2 2 2336 2337 
2 2378 1 2377  
2 2379 1 2377  
0 2380 4 2 2 2338 2339 
2 2381 1 2380  
2 2382 1 2380  
0 2383 4 2 2 2340 2341 
2 2384 1 2383  
2 2385 1 2383  
0 2386 4 2 2 2342 2343 
2 2387 1 2386  
2 2388 1 2386  
0 2389 4 2 2 2344 2345 
2 2390 1 2389  
2 2391 1 2389  
0 2392 4 2 2 2346 2347 
2 2393 1 2392  
2 2394 1 2392  
0 2395 4 2 2 2348 2349 
2 2396 1 2395  
2 2397 1 2395  
0 2398 4 3 2 2351 1132 
2 2399 1 2398  
2 2400 1 2398  
2 2401 1 2398  
0 2402 4 1 2 2321 2354 
0 2403 4 1 2 2355 1181 
0 2404 4 2 2 2220 2356 
2 2405 1 2404  
2 2406 1 2404  
0 2407 4 2 2 2357 2358 
2 2408 1 2407  
2 2409 1 2407  
0 2410 4 3 2 1276 2360 
2 2411 1 2410  
2 2412 1 2410  
2 2413 1 2410  
0 2414 4 3 2 2363 556 
2 2415 1 2414  
2 2416 1 2414  
2 2417 1 2414  
0 2418 4 3 2 2366 604 
2 2419 1 2418  
2 2420 1 2418  
2 2421 1 2418  
0 2422 4 3 2 2369 652 
2 2423 1 2422  
2 2424 1 2422  
2 2425 1 2422  
0 2426 4 3 2 2372 700 
2 2427 1 2426  
2 2428 1 2426  
2 2429 1 2426  
0 2430 4 3 2 2375 748 
2 2431 1 2430  
2 2432 1 2430  
2 2433 1 2430  
0 2434 4 3 2 2378 796 
2 2435 1 2434  
2 2436 1 2434  
2 2437 1 2434  
0 2438 4 3 2 2381 844 
2 2439 1 2438  
2 2440 1 2438  
2 2441 1 2438  
0 2442 4 3 2 2384 892 
2 2443 1 2442  
2 2444 1 2442  
2 2445 1 2442  
0 2446 4 3 2 2387 940 
2 2447 1 2446  
2 2448 1 2446  
2 2449 1 2446  
0 2450 4 3 2 2390 988 
2 2451 1 2450  
2 2452 1 2450  
2 2453 1 2450  
0 2454 4 3 2 2393 1036 
2 2455 1 2454  
2 2456 1 2454  
2 2457 1 2454  
0 2458 4 3 2 2396 1084 
2 2459 1 2458  
2 2460 1 2458  
2 2461 1 2458  
0 2462 4 1 2 2352 2399 
0 2463 4 1 2 2400 1133 
0 2464 4 2 2 2263 2401 
2 2465 1 2464  
2 2466 1 2464  
0 2467 4 2 2 2402 2403 
2 2468 1 2467  
2 2469 1 2467  
0 2470 4 3 2 2408 2405 
2 2471 1 2470  
2 2472 1 2470  
2 2473 1 2470  
0 2474 4 1 2 1277 2411 
0 2475 4 1 2 2412 2361 
0 2476 4 1 2 2364 2415 
0 2477 4 1 2 2416 557 
0 2478 4 2 2 2272 2417 
2 2479 1 2478  
2 2480 1 2478  
0 2481 4 1 2 2367 2419 
0 2482 4 1 2 2420 605 
0 2483 4 2 2 2276 2421 
2 2484 1 2483  
2 2485 1 2483  
0 2486 4 1 2 2370 2423 
0 2487 4 1 2 2424 653 
0 2488 4 2 2 2280 2425 
2 2489 1 2488  
2 2490 1 2488  
0 2491 4 1 2 2373 2427 
0 2492 4 1 2 2428 701 
0 2493 4 2 2 2284 2429 
2 2494 1 2493  
2 2495 1 2493  
0 2496 4 1 2 2376 2431 
0 2497 4 1 2 2432 749 
0 2498 4 2 2 2288 2433 
2 2499 1 2498  
2 2500 1 2498  
0 2501 4 1 2 2379 2435 
0 2502 4 1 2 2436 797 
0 2503 4 2 2 2292 2437 
2 2504 1 2503  
2 2505 1 2503  
0 2506 4 1 2 2382 2439 
0 2507 4 1 2 2440 845 
0 2508 4 2 2 2296 2441 
2 2509 1 2508  
2 2510 1 2508  
0 2511 4 1 2 2385 2443 
0 2512 4 1 2 2444 893 
0 2513 4 2 2 2300 2445 
2 2514 1 2513  
2 2515 1 2513  
0 2516 4 1 2 2388 2447 
0 2517 4 1 2 2448 941 
0 2518 4 2 2 2304 2449 
2 2519 1 2518  
2 2520 1 2518  
0 2521 4 1 2 2391 2451 
0 2522 4 1 2 2452 989 
0 2523 4 2 2 2308 2453 
2 2524 1 2523  
2 2525 1 2523  
0 2526 4 1 2 2394 2455 
0 2527 4 1 2 2456 1037 
0 2528 4 2 2 2312 2457 
2 2529 1 2528  
2 2530 1 2528  
0 2531 4 1 2 2397 2459 
0 2532 4 1 2 2460 1085 
0 2533 4 2 2 2316 2461 
2 2534 1 2533  
2 2535 1 2533  
0 2536 4 2 2 2462 2463 
2 2537 1 2536  
2 2538 1 2536  
0 2539 4 3 2 2468 2465 
2 2540 1 2539  
2 2541 1 2539  
2 2542 1 2539  
0 2543 4 1 2 2409 2471 
0 2544 4 1 2 2472 2406 
0 2545 4 2 2 2474 2475 
2 2546 1 2545  
2 2547 1 2545  
3 2548 4 0 2 2476 2477 
0 2549 4 2 2 2481 2482 
2 2550 1 2549  
2 2551 1 2549  
0 2552 4 2 2 2486 2487 
2 2553 1 2552  
2 2554 1 2552  
0 2555 4 2 2 2491 2492 
2 2556 1 2555  
2 2557 1 2555  
0 2558 4 2 2 2496 2497 
2 2559 1 2558  
2 2560 1 2558  
0 2561 4 2 2 2501 2502 
2 2562 1 2561  
2 2563 1 2561  
0 2564 4 2 2 2506 2507 
2 2565 1 2564  
2 2566 1 2564  
0 2567 4 2 2 2511 2512 
2 2568 1 2567  
2 2569 1 2567  
0 2570 4 2 2 2516 2517 
2 2571 1 2570  
2 2572 1 2570  
0 2573 4 2 2 2521 2522 
2 2574 1 2573  
2 2575 1 2573  
0 2576 4 2 2 2526 2527 
2 2577 1 2576  
2 2578 1 2576  
0 2579 4 2 2 2531 2532 
2 2580 1 2579  
2 2581 1 2579  
0 2582 4 3 2 2537 2534 
2 2583 1 2582  
2 2584 1 2582  
2 2585 1 2582  
0 2586 4 1 2 2469 2540 
0 2587 4 1 2 2541 2466 
0 2588 4 2 2 2543 2544 
2 2589 1 2588  
2 2590 1 2588  
0 2591 4 3 2 2546 1231 
2 2592 1 2591  
2 2593 1 2591  
2 2594 1 2591  
0 2595 4 3 2 2550 2479 
2 2596 1 2595  
2 2597 1 2595  
2 2598 1 2595  
0 2599 4 3 2 2553 2484 
2 2600 1 2599  
2 2601 1 2599  
2 2602 1 2599  
0 2603 4 3 2 2556 2489 
2 2604 1 2603  
2 2605 1 2603  
2 2606 1 2603  
0 2607 4 3 2 2559 2494 
2 2608 1 2607  
2 2609 1 2607  
2 2610 1 2607  
0 2611 4 3 2 2562 2499 
2 2612 1 2611  
2 2613 1 2611  
2 2614 1 2611  
0 2615 4 3 2 2565 2504 
2 2616 1 2615  
2 2617 1 2615  
2 2618 1 2615  
0 2619 4 3 2 2568 2509 
2 2620 1 2619  
2 2621 1 2619  
2 2622 1 2619  
0 2623 4 3 2 2571 2514 
2 2624 1 2623  
2 2625 1 2623  
2 2626 1 2623  
0 2627 4 3 2 2574 2519 
2 2628 1 2627  
2 2629 1 2627  
2 2630 1 2627  
0 2631 4 3 2 2577 2524 
2 2632 1 2631  
2 2633 1 2631  
2 2634 1 2631  
0 2635 4 3 2 2580 2529 
2 2636 1 2635  
2 2637 1 2635  
2 2638 1 2635  
0 2639 4 1 2 2538 2583 
0 2640 4 1 2 2584 2535 
0 2641 4 2 2 2586 2587 
2 2642 1 2641  
2 2643 1 2641  
0 2644 4 3 2 2589 1183 
2 2645 1 2644  
2 2646 1 2644  
2 2647 1 2644  
0 2648 4 1 2 2547 2592 
0 2649 4 1 2 2593 1232 
0 2650 4 2 2 2413 2594 
2 2651 1 2650  
2 2652 1 2650  
0 2653 4 1 2 2551 2596 
0 2654 4 1 2 2597 2480 
0 2655 4 1 2 2554 2600 
0 2656 4 1 2 2601 2485 
0 2657 4 1 2 2557 2604 
0 2658 4 1 2 2605 2490 
0 2659 4 1 2 2560 2608 
0 2660 4 1 2 2609 2495 
0 2661 4 1 2 2563 2612 
0 2662 4 1 2 2613 2500 
0 2663 4 1 2 2566 2616 
0 2664 4 1 2 2617 2505 
0 2665 4 1 2 2569 2620 
0 2666 4 1 2 2621 2510 
0 2667 4 1 2 2572 2624 
0 2668 4 1 2 2625 2515 
0 2669 4 1 2 2575 2628 
0 2670 4 1 2 2629 2520 
0 2671 4 1 2 2578 2632 
0 2672 4 1 2 2633 2525 
0 2673 4 1 2 2581 2636 
0 2674 4 1 2 2637 2530 
0 2675 4 2 2 2639 2640 
2 2676 1 2675  
2 2677 1 2675  
0 2678 4 3 2 2642 1135 
2 2679 1 2678  
2 2680 1 2678  
2 2681 1 2678  
0 2682 4 1 2 2590 2645 
0 2683 4 1 2 2646 1184 
0 2684 4 2 2 2473 2647 
2 2685 1 2684  
2 2686 1 2684  
0 2687 4 2 2 2648 2649 
2 2688 1 2687  
2 2689 1 2687  
0 2690 4 3 2 1279 2651 
2 2691 1 2690  
2 2692 1 2690  
2 2693 1 2690  
0 2694 4 2 2 2653 2654 
2 2695 1 2694  
2 2696 1 2694  
0 2697 4 2 2 2655 2656 
2 2698 1 2697  
2 2699 1 2697  
0 2700 4 2 2 2657 2658 
2 2701 1 2700  
2 2702 1 2700  
0 2703 4 2 2 2659 2660 
2 2704 1 2703  
2 2705 1 2703  
0 2706 4 2 2 2661 2662 
2 2707 1 2706  
2 2708 1 2706  
0 2709 4 2 2 2663 2664 
2 2710 1 2709  
2 2711 1 2709  
0 2712 4 2 2 2665 2666 
2 2713 1 2712  
2 2714 1 2712  
0 2715 4 2 2 2667 2668 
2 2716 1 2715  
2 2717 1 2715  
0 2718 4 2 2 2669 2670 
2 2719 1 2718  
2 2720 1 2718  
0 2721 4 2 2 2671 2672 
2 2722 1 2721  
2 2723 1 2721  
0 2724 4 2 2 2673 2674 
2 2725 1 2724  
2 2726 1 2724  
0 2727 4 3 2 2676 1087 
2 2728 1 2727  
2 2729 1 2727  
2 2730 1 2727  
0 2731 4 1 2 2643 2679 
0 2732 4 1 2 2680 1136 
0 2733 4 2 2 2542 2681 
2 2734 1 2733  
2 2735 1 2733  
0 2736 4 2 2 2682 2683 
2 2737 1 2736  
2 2738 1 2736  
0 2739 4 3 2 2688 2685 
2 2740 1 2739  
2 2741 1 2739  
2 2742 1 2739  
0 2743 4 1 2 1280 2691 
0 2744 4 1 2 2692 2652 
0 2745 4 3 2 2695 559 
2 2746 1 2745  
2 2747 1 2745  
2 2748 1 2745  
0 2749 4 3 2 2698 607 
2 2750 1 2749  
2 2751 1 2749  
2 2752 1 2749  
0 2753 4 3 2 2701 655 
2 2754 1 2753  
2 2755 1 2753  
2 2756 1 2753  
0 2757 4 3 2 2704 703 
2 2758 1 2757  
2 2759 1 2757  
2 2760 1 2757  
0 2761 4 3 2 2707 751 
2 2762 1 2761  
2 2763 1 2761  
2 2764 1 2761  
0 2765 4 3 2 2710 799 
2 2766 1 2765  
2 2767 1 2765  
2 2768 1 2765  
0 2769 4 3 2 2713 847 
2 2770 1 2769  
2 2771 1 2769  
2 2772 1 2769  
0 2773 4 3 2 2716 895 
2 2774 1 2773  
2 2775 1 2773  
2 2776 1 2773  
0 2777 4 3 2 2719 943 
2 2778 1 2777  
2 2779 1 2777  
2 2780 1 2777  
0 2781 4 3 2 2722 991 
2 2782 1 2781  
2 2783 1 2781  
2 2784 1 2781  
0 2785 4 3 2 2725 1039 
2 2786 1 2785  
2 2787 1 2785  
2 2788 1 2785  
0 2789 4 1 2 2677 2728 
0 2790 4 1 2 2729 1088 
0 2791 4 2 2 2585 2730 
2 2792 1 2791  
2 2793 1 2791  
0 2794 4 2 2 2731 2732 
2 2795 1 2794  
2 2796 1 2794  
0 2797 4 3 2 2737 2734 
2 2798 1 2797  
2 2799 1 2797  
2 2800 1 2797  
0 2801 4 1 2 2689 2740 
0 2802 4 1 2 2741 2686 
0 2803 4 2 2 2743 2744 
2 2804 1 2803  
2 2805 1 2803  
0 2806 4 1 2 2696 2746 
0 2807 4 1 2 2747 560 
0 2808 4 2 2 2598 2748 
2 2809 1 2808  
2 2810 1 2808  
0 2811 4 1 2 2699 2750 
0 2812 4 1 2 2751 608 
0 2813 4 2 2 2602 2752 
2 2814 1 2813  
2 2815 1 2813  
0 2816 4 1 2 2702 2754 
0 2817 4 1 2 2755 656 
0 2818 4 2 2 2606 2756 
2 2819 1 2818  
2 2820 1 2818  
0 2821 4 1 2 2705 2758 
0 2822 4 1 2 2759 704 
0 2823 4 2 2 2610 2760 
2 2824 1 2823  
2 2825 1 2823  
0 2826 4 1 2 2708 2762 
0 2827 4 1 2 2763 752 
0 2828 4 2 2 2614 2764 
2 2829 1 2828  
2 2830 1 2828  
0 2831 4 1 2 2711 2766 
0 2832 4 1 2 2767 800 
0 2833 4 2 2 2618 2768 
2 2834 1 2833  
2 2835 1 2833  
0 2836 4 1 2 2714 2770 
0 2837 4 1 2 2771 848 
0 2838 4 2 2 2622 2772 
2 2839 1 2838  
2 2840 1 2838  
0 2841 4 1 2 2717 2774 
0 2842 4 1 2 2775 896 
0 2843 4 2 2 2626 2776 
2 2844 1 2843  
2 2845 1 2843  
0 2846 4 1 2 2720 2778 
0 2847 4 1 2 2779 944 
0 2848 4 2 2 2630 2780 
2 2849 1 2848  
2 2850 1 2848  
0 2851 4 1 2 2723 2782 
0 2852 4 1 2 2783 992 
0 2853 4 2 2 2634 2784 
2 2854 1 2853  
2 2855 1 2853  
0 2856 4 1 2 2726 2786 
0 2857 4 1 2 2787 1040 
0 2858 4 2 2 2638 2788 
2 2859 1 2858  
2 2860 1 2858  
0 2861 4 2 2 2789 2790 
2 2862 1 2861  
2 2863 1 2861  
0 2864 4 3 2 2795 2792 
2 2865 1 2864  
2 2866 1 2864  
2 2867 1 2864  
0 2868 4 1 2 2738 2798 
0 2869 4 1 2 2799 2735 
0 2870 4 2 2 2801 2802 
2 2871 1 2870  
2 2872 1 2870  
0 2873 4 3 2 2804 1234 
2 2874 1 2873  
2 2875 1 2873  
2 2876 1 2873  
3 2877 4 0 2 2806 2807 
0 2878 4 2 2 2811 2812 
2 2879 1 2878  
2 2880 1 2878  
0 2881 4 2 2 2816 2817 
2 2882 1 2881  
2 2883 1 2881  
0 2884 4 2 2 2821 2822 
2 2885 1 2884  
2 2886 1 2884  
0 2887 4 2 2 2826 2827 
2 2888 1 2887  
2 2889 1 2887  
0 2890 4 2 2 2831 2832 
2 2891 1 2890  
2 2892 1 2890  
0 2893 4 2 2 2836 2837 
2 2894 1 2893  
2 2895 1 2893  
0 2896 4 2 2 2841 2842 
2 2897 1 2896  
2 2898 1 2896  
0 2899 4 2 2 2846 2847 
2 2900 1 2899  
2 2901 1 2899  
0 2902 4 2 2 2851 2852 
2 2903 1 2902  
2 2904 1 2902  
0 2905 4 2 2 2856 2857 
2 2906 1 2905  
2 2907 1 2905  
0 2908 4 3 2 2862 2859 
2 2909 1 2908  
2 2910 1 2908  
2 2911 1 2908  
0 2912 4 1 2 2796 2865 
0 2913 4 1 2 2866 2793 
0 2914 4 2 2 2868 2869 
2 2915 1 2914  
2 2916 1 2914  
0 2917 4 3 2 2871 1186 
2 2918 1 2917  
2 2919 1 2917  
2 2920 1 2917  
0 2921 4 1 2 2805 2874 
0 2922 4 1 2 2875 1235 
0 2923 4 2 2 2693 2876 
2 2924 1 2923  
2 2925 1 2923  
0 2926 4 3 2 2879 2809 
2 2927 1 2926  
2 2928 1 2926  
2 2929 1 2926  
0 2930 4 3 2 2882 2814 
2 2931 1 2930  
2 2932 1 2930  
2 2933 1 2930  
0 2934 4 3 2 2885 2819 
2 2935 1 2934  
2 2936 1 2934  
2 2937 1 2934  
0 2938 4 3 2 2888 2824 
2 2939 1 2938  
2 2940 1 2938  
2 2941 1 2938  
0 2942 4 3 2 2891 2829 
2 2943 1 2942  
2 2944 1 2942  
2 2945 1 2942  
0 2946 4 3 2 2894 2834 
2 2947 1 2946  
2 2948 1 2946  
2 2949 1 2946  
0 2950 4 3 2 2897 2839 
2 2951 1 2950  
2 2952 1 2950  
2 2953 1 2950  
0 2954 4 3 2 2900 2844 
2 2955 1 2954  
2 2956 1 2954  
2 2957 1 2954  
0 2958 4 3 2 2903 2849 
2 2959 1 2958  
2 2960 1 2958  
2 2961 1 2958  
0 2962 4 3 2 2906 2854 
2 2963 1 2962  
2 2964 1 2962  
2 2965 1 2962  
0 2966 4 1 2 2863 2909 
0 2967 4 1 2 2910 2860 
0 2968 4 2 2 2912 2913 
2 2969 1 2968  
2 2970 1 2968  
0 2971 4 3 2 2915 1138 
2 2972 1 2971  
2 2973 1 2971  
2 2974 1 2971  
0 2975 4 1 2 2872 2918 
0 2976 4 1 2 2919 1187 
0 2977 4 2 2 2742 2920 
2 2978 1 2977  
2 2979 1 2977  
0 2980 4 2 2 2921 2922 
2 2981 1 2980  
2 2982 1 2980  
0 2983 4 3 2 1282 2924 
2 2984 1 2983  
2 2985 1 2983  
2 2986 1 2983  
0 2987 4 1 2 2880 2927 
0 2988 4 1 2 2928 2810 
0 2989 4 1 2 2883 2931 
0 2990 4 1 2 2932 2815 
0 2991 4 1 2 2886 2935 
0 2992 4 1 2 2936 2820 
0 2993 4 1 2 2889 2939 
0 2994 4 1 2 2940 2825 
0 2995 4 1 2 2892 2943 
0 2996 4 1 2 2944 2830 
0 2997 4 1 2 2895 2947 
0 2998 4 1 2 2948 2835 
0 2999 4 1 2 2898 2951 
0 3000 4 1 2 2952 2840 
0 3001 4 1 2 2901 2955 
0 3002 4 1 2 2956 2845 
0 3003 4 1 2 2904 2959 
0 3004 4 1 2 2960 2850 
0 3005 4 1 2 2907 2963 
0 3006 4 1 2 2964 2855 
0 3007 4 2 2 2966 2967 
2 3008 1 3007  
2 3009 1 3007  
0 3010 4 3 2 2969 1090 
2 3011 1 3010  
2 3012 1 3010  
2 3013 1 3010  
0 3014 4 1 2 2916 2972 
0 3015 4 1 2 2973 1139 
0 3016 4 2 2 2800 2974 
2 3017 1 3016  
2 3018 1 3016  
0 3019 4 2 2 2975 2976 
2 3020 1 3019  
2 3021 1 3019  
0 3022 4 3 2 2981 2978 
2 3023 1 3022  
2 3024 1 3022  
2 3025 1 3022  
0 3026 4 1 2 1283 2984 
0 3027 4 1 2 2985 2925 
0 3028 4 2 2 2987 2988 
2 3029 1 3028  
2 3030 1 3028  
0 3031 4 2 2 2989 2990 
2 3032 1 3031  
2 3033 1 3031  
0 3034 4 2 2 2991 2992 
2 3035 1 3034  
2 3036 1 3034  
0 3037 4 2 2 2993 2994 
2 3038 1 3037  
2 3039 1 3037  
0 3040 4 2 2 2995 2996 
2 3041 1 3040  
2 3042 1 3040  
0 3043 4 2 2 2997 2998 
2 3044 1 3043  
2 3045 1 3043  
0 3046 4 2 2 2999 3000 
2 3047 1 3046  
2 3048 1 3046  
0 3049 4 2 2 3001 3002 
2 3050 1 3049  
2 3051 1 3049  
0 3052 4 2 2 3003 3004 
2 3053 1 3052  
2 3054 1 3052  
0 3055 4 2 2 3005 3006 
2 3056 1 3055  
2 3057 1 3055  
0 3058 4 3 2 3008 1042 
2 3059 1 3058  
2 3060 1 3058  
2 3061 1 3058  
0 3062 4 1 2 2970 3011 
0 3063 4 1 2 3012 1091 
0 3064 4 2 2 2867 3013 
2 3065 1 3064  
2 3066 1 3064  
0 3067 4 2 2 3014 3015 
2 3068 1 3067  
2 3069 1 3067  
0 3070 4 3 2 3020 3017 
2 3071 1 3070  
2 3072 1 3070  
2 3073 1 3070  
0 3074 4 1 2 2982 3023 
0 3075 4 1 2 3024 2979 
0 3076 4 2 2 3026 3027 
2 3077 1 3076  
2 3078 1 3076  
0 3079 4 3 2 3029 562 
2 3080 1 3079  
2 3081 1 3079  
2 3082 1 3079  
0 3083 4 3 2 3032 610 
2 3084 1 3083  
2 3085 1 3083  
2 3086 1 3083  
0 3087 4 3 2 3035 658 
2 3088 1 3087  
2 3089 1 3087  
2 3090 1 3087  
0 3091 4 3 2 3038 706 
2 3092 1 3091  
2 3093 1 3091  
2 3094 1 3091  
0 3095 4 3 2 3041 754 
2 3096 1 3095  
2 3097 1 3095  
2 3098 1 3095  
0 3099 4 3 2 3044 802 
2 3100 1 3099  
2 3101 1 3099  
2 3102 1 3099  
0 3103 4 3 2 3047 850 
2 3104 1 3103  
2 3105 1 3103  
2 3106 1 3103  
0 3107 4 3 2 3050 898 
2 3108 1 3107  
2 3109 1 3107  
2 3110 1 3107  
0 3111 4 3 2 3053 946 
2 3112 1 3111  
2 3113 1 3111  
2 3114 1 3111  
0 3115 4 3 2 3056 994 
2 3116 1 3115  
2 3117 1 3115  
2 3118 1 3115  
0 3119 4 1 2 3009 3059 
0 3120 4 1 2 3060 1043 
0 3121 4 2 2 2911 3061 
2 3122 1 3121  
2 3123 1 3121  
0 3124 4 2 2 3062 3063 
2 3125 1 3124  
2 3126 1 3124  
0 3127 4 3 2 3068 3065 
2 3128 1 3127  
2 3129 1 3127  
2 3130 1 3127  
0 3131 4 1 2 3021 3071 
0 3132 4 1 2 3072 3018 
0 3133 4 2 2 3074 3075 
2 3134 1 3133  
2 3135 1 3133  
0 3136 4 3 2 3077 1237 
2 3137 1 3136  
2 3138 1 3136  
2 3139 1 3136  
0 3140 4 1 2 3030 3080 
0 3141 4 1 2 3081 563 
0 3142 4 2 2 2929 3082 
2 3143 1 3142  
2 3144 1 3142  
0 3145 4 1 2 3033 3084 
0 3146 4 1 2 3085 611 
0 3147 4 2 2 2933 3086 
2 3148 1 3147  
2 3149 1 3147  
0 3150 4 1 2 3036 3088 
0 3151 4 1 2 3089 659 
0 3152 4 2 2 2937 3090 
2 3153 1 3152  
2 3154 1 3152  
0 3155 4 1 2 3039 3092 
0 3156 4 1 2 3093 707 
0 3157 4 2 2 2941 3094 
2 3158 1 3157  
2 3159 1 3157  
0 3160 4 1 2 3042 3096 
0 3161 4 1 2 3097 755 
0 3162 4 2 2 2945 3098 
2 3163 1 3162  
2 3164 1 3162  
0 3165 4 1 2 3045 3100 
0 3166 4 1 2 3101 803 
0 3167 4 2 2 2949 3102 
2 3168 1 3167  
2 3169 1 3167  
0 3170 4 1 2 3048 3104 
0 3171 4 1 2 3105 851 
0 3172 4 2 2 2953 3106 
2 3173 1 3172  
2 3174 1 3172  
0 3175 4 1 2 3051 3108 
0 3176 4 1 2 3109 899 
0 3177 4 2 2 2957 3110 
2 3178 1 3177  
2 3179 1 3177  
0 3180 4 1 2 3054 3112 
0 3181 4 1 2 3113 947 
0 3182 4 2 2 2961 3114 
2 3183 1 3182  
2 3184 1 3182  
0 3185 4 1 2 3057 3116 
0 3186 4 1 2 3117 995 
0 3187 4 2 2 2965 3118 
2 3188 1 3187  
2 3189 1 3187  
0 3190 4 2 2 3119 3120 
2 3191 1 3190  
2 3192 1 3190  
0 3193 4 3 2 3125 3122 
2 3194 1 3193  
2 3195 1 3193  
2 3196 1 3193  
0 3197 4 1 2 3069 3128 
0 3198 4 1 2 3129 3066 
0 3199 4 2 2 3131 3132 
2 3200 1 3199  
2 3201 1 3199  
0 3202 4 3 2 3134 1189 
2 3203 1 3202  
2 3204 1 3202  
2 3205 1 3202  
0 3206 4 1 2 3078 3137 
0 3207 4 1 2 3138 1238 
0 3208 4 2 2 2986 3139 
2 3209 1 3208  
2 3210 1 3208  
3 3211 4 0 2 3140 3141 
0 3212 4 2 2 3145 3146 
2 3213 1 3212  
2 3214 1 3212  
0 3215 4 2 2 3150 3151 
2 3216 1 3215  
2 3217 1 3215  
0 3218 4 2 2 3155 3156 
2 3219 1 3218  
2 3220 1 3218  
0 3221 4 2 2 3160 3161 
2 3222 1 3221  
2 3223 1 3221  
0 3224 4 2 2 3165 3166 
2 3225 1 3224  
2 3226 1 3224  
0 3227 4 2 2 3170 3171 
2 3228 1 3227  
2 3229 1 3227  
0 3230 4 2 2 3175 3176 
2 3231 1 3230  
2 3232 1 3230  
0 3233 4 2 2 3180 3181 
2 3234 1 3233  
2 3235 1 3233  
0 3236 4 2 2 3185 3186 
2 3237 1 3236  
2 3238 1 3236  
0 3239 4 3 2 3191 3188 
2 3240 1 3239  
2 3241 1 3239  
2 3242 1 3239  
0 3243 4 1 2 3126 3194 
0 3244 4 1 2 3195 3123 
0 3245 4 2 2 3197 3198 
2 3246 1 3245  
2 3247 1 3245  
0 3248 4 3 2 3200 1141 
2 3249 1 3248  
2 3250 1 3248  
2 3251 1 3248  
0 3252 4 1 2 3135 3203 
0 3253 4 1 2 3204 1190 
0 3254 4 2 2 3025 3205 
2 3255 1 3254  
2 3256 1 3254  
0 3257 4 2 2 3206 3207 
2 3258 1 3257  
2 3259 1 3257  
0 3260 4 3 2 1285 3209 
2 3261 1 3260  
2 3262 1 3260  
2 3263 1 3260  
0 3264 4 3 2 3213 3143 
2 3265 1 3264  
2 3266 1 3264  
2 3267 1 3264  
0 3268 4 3 2 3216 3148 
2 3269 1 3268  
2 3270 1 3268  
2 3271 1 3268  
0 3272 4 3 2 3219 3153 
2 3273 1 3272  
2 3274 1 3272  
2 3275 1 3272  
0 3276 4 3 2 3222 3158 
2 3277 1 3276  
2 3278 1 3276  
2 3279 1 3276  
0 3280 4 3 2 3225 3163 
2 3281 1 3280  
2 3282 1 3280  
2 3283 1 3280  
0 3284 4 3 2 3228 3168 
2 3285 1 3284  
2 3286 1 3284  
2 3287 1 3284  
0 3288 4 3 2 3231 3173 
2 3289 1 3288  
2 3290 1 3288  
2 3291 1 3288  
0 3292 4 3 2 3234 3178 
2 3293 1 3292  
2 3294 1 3292  
2 3295 1 3292  
0 3296 4 3 2 3237 3183 
2 3297 1 3296  
2 3298 1 3296  
2 3299 1 3296  
0 3300 4 1 2 3192 3240 
0 3301 4 1 2 3241 3189 
0 3302 4 2 2 3243 3244 
2 3303 1 3302  
2 3304 1 3302  
0 3305 4 3 2 3246 1093 
2 3306 1 3305  
2 3307 1 3305  
2 3308 1 3305  
0 3309 4 1 2 3201 3249 
0 3310 4 1 2 3250 1142 
0 3311 4 2 2 3073 3251 
2 3312 1 3311  
2 3313 1 3311  
0 3314 4 2 2 3252 3253 
2 3315 1 3314  
2 3316 1 3314  
0 3317 4 3 2 3258 3255 
2 3318 1 3317  
2 3319 1 3317  
2 3320 1 3317  
0 3321 4 1 2 1286 3261 
0 3322 4 1 2 3262 3210 
0 3323 4 1 2 3214 3265 
0 3324 4 1 2 3266 3144 
0 3325 4 1 2 3217 3269 
0 3326 4 1 2 3270 3149 
0 3327 4 1 2 3220 3273 
0 3328 4 1 2 3274 3154 
0 3329 4 1 2 3223 3277 
0 3330 4 1 2 3278 3159 
0 3331 4 1 2 3226 3281 
0 3332 4 1 2 3282 3164 
0 3333 4 1 2 3229 3285 
0 3334 4 1 2 3286 3169 
0 3335 4 1 2 3232 3289 
0 3336 4 1 2 3290 3174 
0 3337 4 1 2 3235 3293 
0 3338 4 1 2 3294 3179 
0 3339 4 1 2 3238 3297 
0 3340 4 1 2 3298 3184 
0 3341 4 2 2 3300 3301 
2 3342 1 3341  
2 3343 1 3341  
0 3344 4 3 2 3303 1045 
2 3345 1 3344  
2 3346 1 3344  
2 3347 1 3344  
0 3348 4 1 2 3247 3306 
0 3349 4 1 2 3307 1094 
0 3350 4 2 2 3130 3308 
2 3351 1 3350  
2 3352 1 3350  
0 3353 4 2 2 3309 3310 
2 3354 1 3353  
2 3355 1 3353  
0 3356 4 3 2 3315 3312 
2 3357 1 3356  
2 3358 1 3356  
2 3359 1 3356  
0 3360 4 1 2 3259 3318 
0 3361 4 1 2 3319 3256 
0 3362 4 2 2 3321 3322 
2 3363 1 3362  
2 3364 1 3362  
0 3365 4 2 2 3323 3324 
2 3366 1 3365  
2 3367 1 3365  
0 3368 4 2 2 3325 3326 
2 3369 1 3368  
2 3370 1 3368  
0 3371 4 2 2 3327 3328 
2 3372 1 3371  
2 3373 1 3371  
0 3374 4 2 2 3329 3330 
2 3375 1 3374  
2 3376 1 3374  
0 3377 4 2 2 3331 3332 
2 3378 1 3377  
2 3379 1 3377  
0 3380 4 2 2 3333 3334 
2 3381 1 3380  
2 3382 1 3380  
0 3383 4 2 2 3335 3336 
2 3384 1 3383  
2 3385 1 3383  
0 3386 4 2 2 3337 3338 
2 3387 1 3386  
2 3388 1 3386  
0 3389 4 2 2 3339 3340 
2 3390 1 3389  
2 3391 1 3389  
0 3392 4 3 2 3342 997 
2 3393 1 3392  
2 3394 1 3392  
2 3395 1 3392  
0 3396 4 1 2 3304 3345 
0 3397 4 1 2 3346 1046 
0 3398 4 2 2 3196 3347 
2 3399 1 3398  
2 3400 1 3398  
0 3401 4 2 2 3348 3349 
2 3402 1 3401  
2 3403 1 3401  
0 3404 4 3 2 3354 3351 
2 3405 1 3404  
2 3406 1 3404  
2 3407 1 3404  
0 3408 4 1 2 3316 3357 
0 3409 4 1 2 3358 3313 
0 3410 4 2 2 3360 3361 
2 3411 1 3410  
2 3412 1 3410  
0 3413 4 3 2 3363 1240 
2 3414 1 3413  
2 3415 1 3413  
2 3416 1 3413  
0 3417 4 3 2 3366 565 
2 3418 1 3417  
2 3419 1 3417  
2 3420 1 3417  
0 3421 4 3 2 3369 613 
2 3422 1 3421  
2 3423 1 3421  
2 3424 1 3421  
0 3425 4 3 2 3372 661 
2 3426 1 3425  
2 3427 1 3425  
2 3428 1 3425  
0 3429 4 3 2 3375 709 
2 3430 1 3429  
2 3431 1 3429  
2 3432 1 3429  
0 3433 4 3 2 3378 757 
2 3434 1 3433  
2 3435 1 3433  
2 3436 1 3433  
0 3437 4 3 2 3381 805 
2 3438 1 3437  
2 3439 1 3437  
2 3440 1 3437  
0 3441 4 3 2 3384 853 
2 3442 1 3441  
2 3443 1 3441  
2 3444 1 3441  
0 3445 4 3 2 3387 901 
2 3446 1 3445  
2 3447 1 3445  
2 3448 1 3445  
0 3449 4 3 2 3390 949 
2 3450 1 3449  
2 3451 1 3449  
2 3452 1 3449  
0 3453 4 1 2 3343 3393 
0 3454 4 1 2 3394 998 
0 3455 4 2 2 3242 3395 
2 3456 1 3455  
2 3457 1 3455  
0 3458 4 2 2 3396 3397 
2 3459 1 3458  
2 3460 1 3458  
0 3461 4 3 2 3402 3399 
2 3462 1 3461  
2 3463 1 3461  
2 3464 1 3461  
0 3465 4 1 2 3355 3405 
0 3466 4 1 2 3406 3352 
0 3467 4 2 2 3408 3409 
2 3468 1 3467  
2 3469 1 3467  
0 3470 4 3 2 3411 1192 
2 3471 1 3470  
2 3472 1 3470  
2 3473 1 3470  
0 3474 4 1 2 3364 3414 
0 3475 4 1 2 3415 1241 
0 3476 4 2 2 3263 3416 
2 3477 1 3476  
2 3478 1 3476  
0 3479 4 1 2 3367 3418 
0 3480 4 1 2 3419 566 
0 3481 4 2 2 3267 3420 
2 3482 1 3481  
2 3483 1 3481  
0 3484 4 1 2 3370 3422 
0 3485 4 1 2 3423 614 
0 3486 4 2 2 3271 3424 
2 3487 1 3486  
2 3488 1 3486  
0 3489 4 1 2 3373 3426 
0 3490 4 1 2 3427 662 
0 3491 4 2 2 3275 3428 
2 3492 1 3491  
2 3493 1 3491  
0 3494 4 1 2 3376 3430 
0 3495 4 1 2 3431 710 
0 3496 4 2 2 3279 3432 
2 3497 1 3496  
2 3498 1 3496  
0 3499 4 1 2 3379 3434 
0 3500 4 1 2 3435 758 
0 3501 4 2 2 3283 3436 
2 3502 1 3501  
2 3503 1 3501  
0 3504 4 1 2 3382 3438 
0 3505 4 1 2 3439 806 
0 3506 4 2 2 3287 3440 
2 3507 1 3506  
2 3508 1 3506  
0 3509 4 1 2 3385 3442 
0 3510 4 1 2 3443 854 
0 3511 4 2 2 3291 3444 
2 3512 1 3511  
2 3513 1 3511  
0 3514 4 1 2 3388 3446 
0 3515 4 1 2 3447 902 
0 3516 4 2 2 3295 3448 
2 3517 1 3516  
2 3518 1 3516  
0 3519 4 1 2 3391 3450 
0 3520 4 1 2 3451 950 
0 3521 4 2 2 3299 3452 
2 3522 1 3521  
2 3523 1 3521  
0 3524 4 2 2 3453 3454 
2 3525 1 3524  
2 3526 1 3524  
0 3527 4 3 2 3459 3456 
2 3528 1 3527  
2 3529 1 3527  
2 3530 1 3527  
0 3531 4 1 2 3403 3462 
0 3532 4 1 2 3463 3400 
0 3533 4 2 2 3465 3466 
2 3534 1 3533  
2 3535 1 3533  
0 3536 4 3 2 3468 1144 
2 3537 1 3536  
2 3538 1 3536  
2 3539 1 3536  
0 3540 4 1 2 3412 3471 
0 3541 4 1 2 3472 1193 
0 3542 4 2 2 3320 3473 
2 3543 1 3542  
2 3544 1 3542  
0 3545 4 2 2 3474 3475 
2 3546 1 3545  
2 3547 1 3545  
0 3548 4 3 2 1288 3477 
2 3549 1 3548  
2 3550 1 3548  
2 3551 1 3548  
3 3552 4 0 2 3479 3480 
0 3553 4 2 2 3484 3485 
2 3554 1 3553  
2 3555 1 3553  
0 3556 4 2 2 3489 3490 
2 3557 1 3556  
2 3558 1 3556  
0 3559 4 2 2 3494 3495 
2 3560 1 3559  
2 3561 1 3559  
0 3562 4 2 2 3499 3500 
2 3563 1 3562  
2 3564 1 3562  
0 3565 4 2 2 3504 3505 
2 3566 1 3565  
2 3567 1 3565  
0 3568 4 2 2 3509 3510 
2 3569 1 3568  
2 3570 1 3568  
0 3571 4 2 2 3514 3515 
2 3572 1 3571  
2 3573 1 3571  
0 3574 4 2 2 3519 3520 
2 3575 1 3574  
2 3576 1 3574  
0 3577 4 3 2 3525 3522 
2 3578 1 3577  
2 3579 1 3577  
2 3580 1 3577  
0 3581 4 1 2 3460 3528 
0 3582 4 1 2 3529 3457 
0 3583 4 2 2 3531 3532 
2 3584 1 3583  
2 3585 1 3583  
0 3586 4 3 2 3534 1096 
2 3587 1 3586  
2 3588 1 3586  
2 3589 1 3586  
0 3590 4 1 2 3469 3537 
0 3591 4 1 2 3538 1145 
0 3592 4 2 2 3359 3539 
2 3593 1 3592  
2 3594 1 3592  
0 3595 4 2 2 3540 3541 
2 3596 1 3595  
2 3597 1 3595  
0 3598 4 3 2 3546 3543 
2 3599 1 3598  
2 3600 1 3598  
2 3601 1 3598  
0 3602 4 1 2 1289 3549 
0 3603 4 1 2 3550 3478 
0 3604 4 3 2 3554 3482 
2 3605 1 3604  
2 3606 1 3604  
2 3607 1 3604  
0 3608 4 3 2 3557 3487 
2 3609 1 3608  
2 3610 1 3608  
2 3611 1 3608  
0 3612 4 3 2 3560 3492 
2 3613 1 3612  
2 3614 1 3612  
2 3615 1 3612  
0 3616 4 3 2 3563 3497 
2 3617 1 3616  
2 3618 1 3616  
2 3619 1 3616  
0 3620 4 3 2 3566 3502 
2 3621 1 3620  
2 3622 1 3620  
2 3623 1 3620  
0 3624 4 3 2 3569 3507 
2 3625 1 3624  
2 3626 1 3624  
2 3627 1 3624  
0 3628 4 3 2 3572 3512 
2 3629 1 3628  
2 3630 1 3628  
2 3631 1 3628  
0 3632 4 3 2 3575 3517 
2 3633 1 3632  
2 3634 1 3632  
2 3635 1 3632  
0 3636 4 1 2 3526 3578 
0 3637 4 1 2 3579 3523 
0 3638 4 2 2 3581 3582 
2 3639 1 3638  
2 3640 1 3638  
0 3641 4 3 2 3584 1048 
2 3642 1 3641  
2 3643 1 3641  
2 3644 1 3641  
0 3645 4 1 2 3535 3587 
0 3646 4 1 2 3588 1097 
0 3647 4 2 2 3407 3589 
2 3648 1 3647  
2 3649 1 3647  
0 3650 4 2 2 3590 3591 
2 3651 1 3650  
2 3652 1 3650  
0 3653 4 3 2 3596 3593 
2 3654 1 3653  
2 3655 1 3653  
2 3656 1 3653  
0 3657 4 1 2 3547 3599 
0 3658 4 1 2 3600 3544 
0 3659 4 2 2 3602 3603 
2 3660 1 3659  
2 3661 1 3659  
0 3662 4 1 2 3555 3605 
0 3663 4 1 2 3606 3483 
0 3664 4 1 2 3558 3609 
0 3665 4 1 2 3610 3488 
0 3666 4 1 2 3561 3613 
0 3667 4 1 2 3614 3493 
0 3668 4 1 2 3564 3617 
0 3669 4 1 2 3618 3498 
0 3670 4 1 2 3567 3621 
0 3671 4 1 2 3622 3503 
0 3672 4 1 2 3570 3625 
0 3673 4 1 2 3626 3508 
0 3674 4 1 2 3573 3629 
0 3675 4 1 2 3630 3513 
0 3676 4 1 2 3576 3633 
0 3677 4 1 2 3634 3518 
0 3678 4 2 2 3636 3637 
2 3679 1 3678  
2 3680 1 3678  
0 3681 4 3 2 3639 1000 
2 3682 1 3681  
2 3683 1 3681  
2 3684 1 3681  
0 3685 4 1 2 3585 3642 
0 3686 4 1 2 3643 1049 
0 3687 4 2 2 3464 3644 
2 3688 1 3687  
2 3689 1 3687  
0 3690 4 2 2 3645 3646 
2 3691 1 3690  
2 3692 1 3690  
0 3693 4 3 2 3651 3648 
2 3694 1 3693  
2 3695 1 3693  
2 3696 1 3693  
0 3697 4 1 2 3597 3654 
0 3698 4 1 2 3655 3594 
0 3699 4 2 2 3657 3658 
2 3700 1 3699  
2 3701 1 3699  
0 3702 4 3 2 3660 1243 
2 3703 1 3702  
2 3704 1 3702  
2 3705 1 3702  
0 3706 4 2 2 3662 3663 
2 3707 1 3706  
2 3708 1 3706  
0 3709 4 2 2 3664 3665 
2 3710 1 3709  
2 3711 1 3709  
0 3712 4 2 2 3666 3667 
2 3713 1 3712  
2 3714 1 3712  
0 3715 4 2 2 3668 3669 
2 3716 1 3715  
2 3717 1 3715  
0 3718 4 2 2 3670 3671 
2 3719 1 3718  
2 3720 1 3718  
0 3721 4 2 2 3672 3673 
2 3722 1 3721  
2 3723 1 3721  
0 3724 4 2 2 3674 3675 
2 3725 1 3724  
2 3726 1 3724  
0 3727 4 2 2 3676 3677 
2 3728 1 3727  
2 3729 1 3727  
0 3730 4 3 2 3679 952 
2 3731 1 3730  
2 3732 1 3730  
2 3733 1 3730  
0 3734 4 1 2 3640 3682 
0 3735 4 1 2 3683 1001 
0 3736 4 2 2 3530 3684 
2 3737 1 3736  
2 3738 1 3736  
0 3739 4 2 2 3685 3686 
2 3740 1 3739  
2 3741 1 3739  
0 3742 4 3 2 3691 3688 
2 3743 1 3742  
2 3744 1 3742  
2 3745 1 3742  
0 3746 4 1 2 3652 3694 
0 3747 4 1 2 3695 3649 
0 3748 4 2 2 3697 3698 
2 3749 1 3748  
2 3750 1 3748  
0 3751 4 3 2 3700 1195 
2 3752 1 3751  
2 3753 1 3751  
2 3754 1 3751  
0 3755 4 1 2 3661 3703 
0 3756 4 1 2 3704 1244 
0 3757 4 2 2 3551 3705 
2 3758 1 3757  
2 3759 1 3757  
0 3760 4 3 2 3707 568 
2 3761 1 3760  
2 3762 1 3760  
2 3763 1 3760  
0 3764 4 3 2 3710 616 
2 3765 1 3764  
2 3766 1 3764  
2 3767 1 3764  
0 3768 4 3 2 3713 664 
2 3769 1 3768  
2 3770 1 3768  
2 3771 1 3768  
0 3772 4 3 2 3716 712 
2 3773 1 3772  
2 3774 1 3772  
2 3775 1 3772  
0 3776 4 3 2 3719 760 
2 3777 1 3776  
2 3778 1 3776  
2 3779 1 3776  
0 3780 4 3 2 3722 808 
2 3781 1 3780  
2 3782 1 3780  
2 3783 1 3780  
0 3784 4 3 2 3725 856 
2 3785 1 3784  
2 3786 1 3784  
2 3787 1 3784  
0 3788 4 3 2 3728 904 
2 3789 1 3788  
2 3790 1 3788  
2 3791 1 3788  
0 3792 4 1 2 3680 3731 
0 3793 4 1 2 3732 953 
0 3794 4 2 2 3580 3733 
2 3795 1 3794  
2 3796 1 3794  
0 3797 4 2 2 3734 3735 
2 3798 1 3797  
2 3799 1 3797  
0 3800 4 3 2 3740 3737 
2 3801 1 3800  
2 3802 1 3800  
2 3803 1 3800  
0 3804 4 1 2 3692 3743 
0 3805 4 1 2 3744 3689 
0 3806 4 2 2 3746 3747 
2 3807 1 3806  
2 3808 1 3806  
0 3809 4 3 2 3749 1147 
2 3810 1 3809  
2 3811 1 3809  
2 3812 1 3809  
0 3813 4 1 2 3701 3752 
0 3814 4 1 2 3753 1196 
0 3815 4 2 2 3601 3754 
2 3816 1 3815  
2 3817 1 3815  
0 3818 4 2 2 3755 3756 
2 3819 1 3818  
2 3820 1 3818  
0 3821 4 3 2 1291 3758 
2 3822 1 3821  
2 3823 1 3821  
2 3824 1 3821  
0 3825 4 1 2 3708 3761 
0 3826 4 1 2 3762 569 
0 3827 4 2 2 3607 3763 
2 3828 1 3827  
2 3829 1 3827  
0 3830 4 1 2 3711 3765 
0 3831 4 1 2 3766 617 
0 3832 4 2 2 3611 3767 
2 3833 1 3832  
2 3834 1 3832  
0 3835 4 1 2 3714 3769 
0 3836 4 1 2 3770 665 
0 3837 4 2 2 3615 3771 
2 3838 1 3837  
2 3839 1 3837  
0 3840 4 1 2 3717 3773 
0 3841 4 1 2 3774 713 
0 3842 4 2 2 3619 3775 
2 3843 1 3842  
2 3844 1 3842  
0 3845 4 1 2 3720 3777 
0 3846 4 1 2 3778 761 
0 3847 4 2 2 3623 3779 
2 3848 1 3847  
2 3849 1 3847  
0 3850 4 1 2 3723 3781 
0 3851 4 1 2 3782 809 
0 3852 4 2 2 3627 3783 
2 3853 1 3852  
2 3854 1 3852  
0 3855 4 1 2 3726 3785 
0 3856 4 1 2 3786 857 
0 3857 4 2 2 3631 3787 
2 3858 1 3857  
2 3859 1 3857  
0 3860 4 1 2 3729 3789 
0 3861 4 1 2 3790 905 
0 3862 4 2 2 3635 3791 
2 3863 1 3862  
2 3864 1 3862  
0 3865 4 2 2 3792 3793 
2 3866 1 3865  
2 3867 1 3865  
0 3868 4 3 2 3798 3795 
2 3869 1 3868  
2 3870 1 3868  
2 3871 1 3868  
0 3872 4 1 2 3741 3801 
0 3873 4 1 2 3802 3738 
0 3874 4 2 2 3804 3805 
2 3875 1 3874  
2 3876 1 3874  
0 3877 4 3 2 3807 1099 
2 3878 1 3877  
2 3879 1 3877  
2 3880 1 3877  
0 3881 4 1 2 3750 3810 
0 3882 4 1 2 3811 1148 
0 3883 4 2 2 3656 3812 
2 3884 1 3883  
2 3885 1 3883  
0 3886 4 2 2 3813 3814 
2 3887 1 3886  
2 3888 1 3886  
0 3889 4 3 2 3819 3816 
2 3890 1 3889  
2 3891 1 3889  
2 3892 1 3889  
0 3893 4 1 2 1292 3822 
0 3894 4 1 2 3823 3759 
3 3895 4 0 2 3825 3826 
0 3896 4 2 2 3830 3831 
2 3897 1 3896  
2 3898 1 3896  
0 3899 4 2 2 3835 3836 
2 3900 1 3899  
2 3901 1 3899  
0 3902 4 2 2 3840 3841 
2 3903 1 3902  
2 3904 1 3902  
0 3905 4 2 2 3845 3846 
2 3906 1 3905  
2 3907 1 3905  
0 3908 4 2 2 3850 3851 
2 3909 1 3908  
2 3910 1 3908  
0 3911 4 2 2 3855 3856 
2 3912 1 3911  
2 3913 1 3911  
0 3914 4 2 2 3860 3861 
2 3915 1 3914  
2 3916 1 3914  
0 3917 4 3 2 3866 3863 
2 3918 1 3917  
2 3919 1 3917  
2 3920 1 3917  
0 3921 4 1 2 3799 3869 
0 3922 4 1 2 3870 3796 
0 3923 4 2 2 3872 3873 
2 3924 1 3923  
2 3925 1 3923  
0 3926 4 3 2 3875 1051 
2 3927 1 3926  
2 3928 1 3926  
2 3929 1 3926  
0 3930 4 1 2 3808 3878 
0 3931 4 1 2 3879 1100 
0 3932 4 2 2 3696 3880 
2 3933 1 3932  
2 3934 1 3932  
0 3935 4 2 2 3881 3882 
2 3936 1 3935  
2 3937 1 3935  
0 3938 4 3 2 3887 3884 
2 3939 1 3938  
2 3940 1 3938  
2 3941 1 3938  
0 3942 4 1 2 3820 3890 
0 3943 4 1 2 3891 3817 
0 3944 4 2 2 3893 3894 
2 3945 1 3944  
2 3946 1 3944  
0 3947 4 3 2 3897 3828 
2 3948 1 3947  
2 3949 1 3947  
2 3950 1 3947  
0 3951 4 3 2 3900 3833 
2 3952 1 3951  
2 3953 1 3951  
2 3954 1 3951  
0 3955 4 3 2 3903 3838 
2 3956 1 3955  
2 3957 1 3955  
2 3958 1 3955  
0 3959 4 3 2 3906 3843 
2 3960 1 3959  
2 3961 1 3959  
2 3962 1 3959  
0 3963 4 3 2 3909 3848 
2 3964 1 3963  
2 3965 1 3963  
2 3966 1 3963  
0 3967 4 3 2 3912 3853 
2 3968 1 3967  
2 3969 1 3967  
2 3970 1 3967  
0 3971 4 3 2 3915 3858 
2 3972 1 3971  
2 3973 1 3971  
2 3974 1 3971  
0 3975 4 1 2 3867 3918 
0 3976 4 1 2 3919 3864 
0 3977 4 2 2 3921 3922 
2 3978 1 3977  
2 3979 1 3977  
0 3980 4 3 2 3924 1003 
2 3981 1 3980  
2 3982 1 3980  
2 3983 1 3980  
0 3984 4 1 2 3876 3927 
0 3985 4 1 2 3928 1052 
0 3986 4 2 2 3745 3929 
2 3987 1 3986  
2 3988 1 3986  
0 3989 4 2 2 3930 3931 
2 3990 1 3989  
2 3991 1 3989  
0 3992 4 3 2 3936 3933 
2 3993 1 3992  
2 3994 1 3992  
2 3995 1 3992  
0 3996 4 1 2 3888 3939 
0 3997 4 1 2 3940 3885 
0 3998 4 2 2 3942 3943 
2 3999 1 3998  
2 4000 1 3998  
0 4001 4 3 2 3945 1246 
2 4002 1 4001  
2 4003 1 4001  
2 4004 1 4001  
0 4005 4 1 2 3898 3948 
0 4006 4 1 2 3949 3829 
0 4007 4 1 2 3901 3952 
0 4008 4 1 2 3953 3834 
0 4009 4 1 2 3904 3956 
0 4010 4 1 2 3957 3839 
0 4011 4 1 2 3907 3960 
0 4012 4 1 2 3961 3844 
0 4013 4 1 2 3910 3964 
0 4014 4 1 2 3965 3849 
0 4015 4 1 2 3913 3968 
0 4016 4 1 2 3969 3854 
0 4017 4 1 2 3916 3972 
0 4018 4 1 2 3973 3859 
0 4019 4 2 2 3975 3976 
2 4020 1 4019  
2 4021 1 4019  
0 4022 4 3 2 3978 955 
2 4023 1 4022  
2 4024 1 4022  
2 4025 1 4022  
0 4026 4 1 2 3925 3981 
0 4027 4 1 2 3982 1004 
0 4028 4 2 2 3803 3983 
2 4029 1 4028  
2 4030 1 4028  
0 4031 4 2 2 3984 3985 
2 4032 1 4031  
2 4033 1 4031  
0 4034 4 3 2 3990 3987 
2 4035 1 4034  
2 4036 1 4034  
2 4037 1 4034  
0 4038 4 1 2 3937 3993 
0 4039 4 1 2 3994 3934 
0 4040 4 2 2 3996 3997 
2 4041 1 4040  
2 4042 1 4040  
0 4043 4 3 2 3999 1198 
2 4044 1 4043  
2 4045 1 4043  
2 4046 1 4043  
0 4047 4 1 2 3946 4002 
0 4048 4 1 2 4003 1247 
0 4049 4 2 2 3824 4004 
2 4050 1 4049  
2 4051 1 4049  
0 4052 4 2 2 4005 4006 
2 4053 1 4052  
2 4054 1 4052  
0 4055 4 2 2 4007 4008 
2 4056 1 4055  
2 4057 1 4055  
0 4058 4 2 2 4009 4010 
2 4059 1 4058  
2 4060 1 4058  
0 4061 4 2 2 4011 4012 
2 4062 1 4061  
2 4063 1 4061  
0 4064 4 2 2 4013 4014 
2 4065 1 4064  
2 4066 1 4064  
0 4067 4 2 2 4015 4016 
2 4068 1 4067  
2 4069 1 4067  
0 4070 4 2 2 4017 4018 
2 4071 1 4070  
2 4072 1 4070  
0 4073 4 3 2 4020 907 
2 4074 1 4073  
2 4075 1 4073  
2 4076 1 4073  
0 4077 4 1 2 3979 4023 
0 4078 4 1 2 4024 956 
0 4079 4 2 2 3871 4025 
2 4080 1 4079  
2 4081 1 4079  
0 4082 4 2 2 4026 4027 
2 4083 1 4082  
2 4084 1 4082  
0 4085 4 3 2 4032 4029 
2 4086 1 4085  
2 4087 1 4085  
2 4088 1 4085  
0 4089 4 1 2 3991 4035 
0 4090 4 1 2 4036 3988 
0 4091 4 2 2 4038 4039 
2 4092 1 4091  
2 4093 1 4091  
0 4094 4 3 2 4041 1150 
2 4095 1 4094  
2 4096 1 4094  
2 4097 1 4094  
0 4098 4 1 2 4000 4044 
0 4099 4 1 2 4045 1199 
0 4100 4 2 2 3892 4046 
2 4101 1 4100  
2 4102 1 4100  
0 4103 4 2 2 4047 4048 
2 4104 1 4103  
2 4105 1 4103  
0 4106 4 3 2 1294 4050 
2 4107 1 4106  
2 4108 1 4106  
2 4109 1 4106  
0 4110 4 3 2 4053 571 
2 4111 1 4110  
2 4112 1 4110  
2 4113 1 4110  
0 4114 4 3 2 4056 619 
2 4115 1 4114  
2 4116 1 4114  
2 4117 1 4114  
0 4118 4 3 2 4059 667 
2 4119 1 4118  
2 4120 1 4118  
2 4121 1 4118  
0 4122 4 3 2 4062 715 
2 4123 1 4122  
2 4124 1 4122  
2 4125 1 4122  
0 4126 4 3 2 4065 763 
2 4127 1 4126  
2 4128 1 4126  
2 4129 1 4126  
0 4130 4 3 2 4068 811 
2 4131 1 4130  
2 4132 1 4130  
2 4133 1 4130  
0 4134 4 3 2 4071 859 
2 4135 1 4134  
2 4136 1 4134  
2 4137 1 4134  
0 4138 4 1 2 4021 4074 
0 4139 4 1 2 4075 908 
0 4140 4 2 2 3920 4076 
2 4141 1 4140  
2 4142 1 4140  
0 4143 4 2 2 4077 4078 
2 4144 1 4143  
2 4145 1 4143  
0 4146 4 3 2 4083 4080 
2 4147 1 4146  
2 4148 1 4146  
2 4149 1 4146  
0 4150 4 1 2 4033 4086 
0 4151 4 1 2 4087 4030 
0 4152 4 2 2 4089 4090 
2 4153 1 4152  
2 4154 1 4152  
0 4155 4 3 2 4092 1102 
2 4156 1 4155  
2 4157 1 4155  
2 4158 1 4155  
0 4159 4 1 2 4042 4095 
0 4160 4 1 2 4096 1151 
0 4161 4 2 2 3941 4097 
2 4162 1 4161  
2 4163 1 4161  
0 4164 4 2 2 4098 4099 
2 4165 1 4164  
2 4166 1 4164  
0 4167 4 3 2 4104 4101 
2 4168 1 4167  
2 4169 1 4167  
2 4170 1 4167  
0 4171 4 1 2 1295 4107 
0 4172 4 1 2 4108 4051 
0 4173 4 1 2 4054 4111 
0 4174 4 1 2 4112 572 
0 4175 4 2 2 3950 4113 
2 4176 1 4175  
2 4177 1 4175  
0 4178 4 1 2 4057 4115 
0 4179 4 1 2 4116 620 
0 4180 4 2 2 3954 4117 
2 4181 1 4180  
2 4182 1 4180  
0 4183 4 1 2 4060 4119 
0 4184 4 1 2 4120 668 
0 4185 4 2 2 3958 4121 
2 4186 1 4185  
2 4187 1 4185  
0 4188 4 1 2 4063 4123 
0 4189 4 1 2 4124 716 
0 4190 4 2 2 3962 4125 
2 4191 1 4190  
2 4192 1 4190  
0 4193 4 1 2 4066 4127 
0 4194 4 1 2 4128 764 
0 4195 4 2 2 3966 4129 
2 4196 1 4195  
2 4197 1 4195  
0 4198 4 1 2 4069 4131 
0 4199 4 1 2 4132 812 
0 4200 4 2 2 3970 4133 
2 4201 1 4200  
2 4202 1 4200  
0 4203 4 1 2 4072 4135 
0 4204 4 1 2 4136 860 
0 4205 4 2 2 3974 4137 
2 4206 1 4205  
2 4207 1 4205  
0 4208 4 2 2 4138 4139 
2 4209 1 4208  
2 4210 1 4208  
0 4211 4 3 2 4144 4141 
2 4212 1 4211  
2 4213 1 4211  
2 4214 1 4211  
0 4215 4 1 2 4084 4147 
0 4216 4 1 2 4148 4081 
0 4217 4 2 2 4150 4151 
2 4218 1 4217  
2 4219 1 4217  
0 4220 4 3 2 4153 1054 
2 4221 1 4220  
2 4222 1 4220  
2 4223 1 4220  
0 4224 4 1 2 4093 4156 
0 4225 4 1 2 4157 1103 
0 4226 4 2 2 3995 4158 
2 4227 1 4226  
2 4228 1 4226  
0 4229 4 2 2 4159 4160 
2 4230 1 4229  
2 4231 1 4229  
0 4232 4 3 2 4165 4162 
2 4233 1 4232  
2 4234 1 4232  
2 4235 1 4232  
0 4236 4 1 2 4105 4168 
0 4237 4 1 2 4169 4102 
0 4238 4 2 2 4171 4172 
2 4239 1 4238  
2 4240 1 4238  
3 4241 4 0 2 4173 4174 
0 4242 4 2 2 4178 4179 
2 4243 1 4242  
2 4244 1 4242  
0 4245 4 2 2 4183 4184 
2 4246 1 4245  
2 4247 1 4245  
0 4248 4 2 2 4188 4189 
2 4249 1 4248  
2 4250 1 4248  
0 4251 4 2 2 4193 4194 
2 4252 1 4251  
2 4253 1 4251  
0 4254 4 2 2 4198 4199 
2 4255 1 4254  
2 4256 1 4254  
0 4257 4 2 2 4203 4204 
2 4258 1 4257  
2 4259 1 4257  
0 4260 4 3 2 4209 4206 
2 4261 1 4260  
2 4262 1 4260  
2 4263 1 4260  
0 4264 4 1 2 4145 4212 
0 4265 4 1 2 4213 4142 
0 4266 4 2 2 4215 4216 
2 4267 1 4266  
2 4268 1 4266  
0 4269 4 3 2 4218 1006 
2 4270 1 4269  
2 4271 1 4269  
2 4272 1 4269  
0 4273 4 1 2 4154 4221 
0 4274 4 1 2 4222 1055 
0 4275 4 2 2 4037 4223 
2 4276 1 4275  
2 4277 1 4275  
0 4278 4 2 2 4224 4225 
2 4279 1 4278  
2 4280 1 4278  
0 4281 4 3 2 4230 4227 
2 4282 1 4281  
2 4283 1 4281  
2 4284 1 4281  
0 4285 4 1 2 4166 4233 
0 4286 4 1 2 4234 4163 
0 4287 4 2 2 4236 4237 
2 4288 1 4287  
2 4289 1 4287  
0 4290 4 3 2 4239 1249 
2 4291 1 4290  
2 4292 1 4290  
2 4293 1 4290  
0 4294 4 3 2 4243 4176 
2 4295 1 4294  
2 4296 1 4294  
2 4297 1 4294  
0 4298 4 3 2 4246 4181 
2 4299 1 4298  
2 4300 1 4298  
2 4301 1 4298  
0 4302 4 3 2 4249 4186 
2 4303 1 4302  
2 4304 1 4302  
2 4305 1 4302  
0 4306 4 3 2 4252 4191 
2 4307 1 4306  
2 4308 1 4306  
2 4309 1 4306  
0 4310 4 3 2 4255 4196 
2 4311 1 4310  
2 4312 1 4310  
2 4313 1 4310  
0 4314 4 3 2 4258 4201 
2 4315 1 4314  
2 4316 1 4314  
2 4317 1 4314  
0 4318 4 1 2 4210 4261 
0 4319 4 1 2 4262 4207 
0 4320 4 2 2 4264 4265 
2 4321 1 4320  
2 4322 1 4320  
0 4323 4 3 2 4267 958 
2 4324 1 4323  
2 4325 1 4323  
2 4326 1 4323  
0 4327 4 1 2 4219 4270 
0 4328 4 1 2 4271 1007 
0 4329 4 2 2 4088 4272 
2 4330 1 4329  
2 4331 1 4329  
0 4332 4 2 2 4273 4274 
2 4333 1 4332  
2 4334 1 4332  
0 4335 4 3 2 4279 4276 
2 4336 1 4335  
2 4337 1 4335  
2 4338 1 4335  
0 4339 4 1 2 4231 4282 
0 4340 4 1 2 4283 4228 
0 4341 4 2 2 4285 4286 
2 4342 1 4341  
2 4343 1 4341  
0 4344 4 3 2 4288 1201 
2 4345 1 4344  
2 4346 1 4344  
2 4347 1 4344  
0 4348 4 1 2 4240 4291 
0 4349 4 1 2 4292 1250 
0 4350 4 2 2 4109 4293 
2 4351 1 4350  
2 4352 1 4350  
0 4353 4 1 2 4244 4295 
0 4354 4 1 2 4296 4177 
0 4355 4 1 2 4247 4299 
0 4356 4 1 2 4300 4182 
0 4357 4 1 2 4250 4303 
0 4358 4 1 2 4304 4187 
0 4359 4 1 2 4253 4307 
0 4360 4 1 2 4308 4192 
0 4361 4 1 2 4256 4311 
0 4362 4 1 2 4312 4197 
0 4363 4 1 2 4259 4315 
0 4364 4 1 2 4316 4202 
0 4365 4 2 2 4318 4319 
2 4366 1 4365  
2 4367 1 4365  
0 4368 4 3 2 4321 910 
2 4369 1 4368  
2 4370 1 4368  
2 4371 1 4368  
0 4372 4 1 2 4268 4324 
0 4373 4 1 2 4325 959 
0 4374 4 2 2 4149 4326 
2 4375 1 4374  
2 4376 1 4374  
0 4377 4 2 2 4327 4328 
2 4378 1 4377  
2 4379 1 4377  
0 4380 4 3 2 4333 4330 
2 4381 1 4380  
2 4382 1 4380  
2 4383 1 4380  
0 4384 4 1 2 4280 4336 
0 4385 4 1 2 4337 4277 
0 4386 4 2 2 4339 4340 
2 4387 1 4386  
2 4388 1 4386  
0 4389 4 3 2 4342 1153 
2 4390 1 4389  
2 4391 1 4389  
2 4392 1 4389  
0 4393 4 1 2 4289 4345 
0 4394 4 1 2 4346 1202 
0 4395 4 2 2 4170 4347 
2 4396 1 4395  
2 4397 1 4395  
0 4398 4 2 2 4348 4349 
2 4399 1 4398  
2 4400 1 4398  
0 4401 4 3 2 1297 4351 
2 4402 1 4401  
2 4403 1 4401  
2 4404 1 4401  
0 4405 4 2 2 4353 4354 
2 4406 1 4405  
2 4407 1 4405  
0 4408 4 2 2 4355 4356 
2 4409 1 4408  
2 4410 1 4408  
0 4411 4 2 2 4357 4358 
2 4412 1 4411  
2 4413 1 4411  
0 4414 4 2 2 4359 4360 
2 4415 1 4414  
2 4416 1 4414  
0 4417 4 2 2 4361 4362 
2 4418 1 4417  
2 4419 1 4417  
0 4420 4 2 2 4363 4364 
2 4421 1 4420  
2 4422 1 4420  
0 4423 4 3 2 4366 862 
2 4424 1 4423  
2 4425 1 4423  
2 4426 1 4423  
0 4427 4 1 2 4322 4369 
0 4428 4 1 2 4370 911 
0 4429 4 2 2 4214 4371 
2 4430 1 4429  
2 4431 1 4429  
0 4432 4 2 2 4372 4373 
2 4433 1 4432  
2 4434 1 4432  
0 4435 4 3 2 4378 4375 
2 4436 1 4435  
2 4437 1 4435  
2 4438 1 4435  
0 4439 4 1 2 4334 4381 
0 4440 4 1 2 4382 4331 
0 4441 4 2 2 4384 4385 
2 4442 1 4441  
2 4443 1 4441  
0 4444 4 3 2 4387 1105 
2 4445 1 4444  
2 4446 1 4444  
2 4447 1 4444  
0 4448 4 1 2 4343 4390 
0 4449 4 1 2 4391 1154 
0 4450 4 2 2 4235 4392 
2 4451 1 4450  
2 4452 1 4450  
0 4453 4 2 2 4393 4394 
2 4454 1 4453  
2 4455 1 4453  
0 4456 4 3 2 4399 4396 
2 4457 1 4456  
2 4458 1 4456  
2 4459 1 4456  
0 4460 4 1 2 1298 4402 
0 4461 4 1 2 4403 4352 
0 4462 4 3 2 4406 574 
2 4463 1 4462  
2 4464 1 4462  
2 4465 1 4462  
0 4466 4 3 2 4409 622 
2 4467 1 4466  
2 4468 1 4466  
2 4469 1 4466  
0 4470 4 3 2 4412 670 
2 4471 1 4470  
2 4472 1 4470  
2 4473 1 4470  
0 4474 4 3 2 4415 718 
2 4475 1 4474  
2 4476 1 4474  
2 4477 1 4474  
0 4478 4 3 2 4418 766 
2 4479 1 4478  
2 4480 1 4478  
2 4481 1 4478  
0 4482 4 3 2 4421 814 
2 4483 1 4482  
2 4484 1 4482  
2 4485 1 4482  
0 4486 4 1 2 4367 4424 
0 4487 4 1 2 4425 863 
0 4488 4 2 2 4263 4426 
2 4489 1 4488  
2 4490 1 4488  
0 4491 4 2 2 4427 4428 
2 4492 1 4491  
2 4493 1 4491  
0 4494 4 3 2 4433 4430 
2 4495 1 4494  
2 4496 1 4494  
2 4497 1 4494  
0 4498 4 1 2 4379 4436 
0 4499 4 1 2 4437 4376 
0 4500 4 2 2 4439 4440 
2 4501 1 4500  
2 4502 1 4500  
0 4503 4 3 2 4442 1057 
2 4504 1 4503  
2 4505 1 4503  
2 4506 1 4503  
0 4507 4 1 2 4388 4445 
0 4508 4 1 2 4446 1106 
0 4509 4 2 2 4284 4447 
2 4510 1 4509  
2 4511 1 4509  
0 4512 4 2 2 4448 4449 
2 4513 1 4512  
2 4514 1 4512  
0 4515 4 3 2 4454 4451 
2 4516 1 4515  
2 4517 1 4515  
2 4518 1 4515  
0 4519 4 1 2 4400 4457 
0 4520 4 1 2 4458 4397 
0 4521 4 2 2 4460 4461 
2 4522 1 4521  
2 4523 1 4521  
0 4524 4 1 2 4407 4463 
0 4525 4 1 2 4464 575 
0 4526 4 2 2 4297 4465 
2 4527 1 4526  
2 4528 1 4526  
0 4529 4 1 2 4410 4467 
0 4530 4 1 2 4468 623 
0 4531 4 2 2 4301 4469 
2 4532 1 4531  
2 4533 1 4531  
0 4534 4 1 2 4413 4471 
0 4535 4 1 2 4472 671 
0 4536 4 2 2 4305 4473 
2 4537 1 4536  
2 4538 1 4536  
0 4539 4 1 2 4416 4475 
0 4540 4 1 2 4476 719 
0 4541 4 2 2 4309 4477 
2 4542 1 4541  
2 4543 1 4541  
0 4544 4 1 2 4419 4479 
0 4545 4 1 2 4480 767 
0 4546 4 2 2 4313 4481 
2 4547 1 4546  
2 4548 1 4546  
0 4549 4 1 2 4422 4483 
0 4550 4 1 2 4484 815 
0 4551 4 2 2 4317 4485 
2 4552 1 4551  
2 4553 1 4551  
0 4554 4 2 2 4486 4487 
2 4555 1 4554  
2 4556 1 4554  
0 4557 4 3 2 4492 4489 
2 4558 1 4557  
2 4559 1 4557  
2 4560 1 4557  
0 4561 4 1 2 4434 4495 
0 4562 4 1 2 4496 4431 
0 4563 4 2 2 4498 4499 
2 4564 1 4563  
2 4565 1 4563  
0 4566 4 3 2 4501 1009 
2 4567 1 4566  
2 4568 1 4566  
2 4569 1 4566  
0 4570 4 1 2 4443 4504 
0 4571 4 1 2 4505 1058 
0 4572 4 2 2 4338 4506 
2 4573 1 4572  
2 4574 1 4572  
0 4575 4 2 2 4507 4508 
2 4576 1 4575  
2 4577 1 4575  
0 4578 4 3 2 4513 4510 
2 4579 1 4578  
2 4580 1 4578  
2 4581 1 4578  
0 4582 4 1 2 4455 4516 
0 4583 4 1 2 4517 4452 
0 4584 4 2 2 4519 4520 
2 4585 1 4584  
2 4586 1 4584  
0 4587 4 3 2 4522 1252 
2 4588 1 4587  
2 4589 1 4587  
2 4590 1 4587  
3 4591 4 0 2 4524 4525 
0 4592 4 2 2 4529 4530 
2 4593 1 4592  
2 4594 1 4592  
0 4595 4 2 2 4534 4535 
2 4596 1 4595  
2 4597 1 4595  
0 4598 4 2 2 4539 4540 
2 4599 1 4598  
2 4600 1 4598  
0 4601 4 2 2 4544 4545 
2 4602 1 4601  
2 4603 1 4601  
0 4604 4 2 2 4549 4550 
2 4605 1 4604  
2 4606 1 4604  
0 4607 4 3 2 4555 4552 
2 4608 1 4607  
2 4609 1 4607  
2 4610 1 4607  
0 4611 4 1 2 4493 4558 
0 4612 4 1 2 4559 4490 
0 4613 4 2 2 4561 4562 
2 4614 1 4613  
2 4615 1 4613  
0 4616 4 3 2 4564 961 
2 4617 1 4616  
2 4618 1 4616  
2 4619 1 4616  
0 4620 4 1 2 4502 4567 
0 4621 4 1 2 4568 1010 
0 4622 4 2 2 4383 4569 
2 4623 1 4622  
2 4624 1 4622  
0 4625 4 2 2 4570 4571 
2 4626 1 4625  
2 4627 1 4625  
0 4628 4 3 2 4576 4573 
2 4629 1 4628  
2 4630 1 4628  
2 4631 1 4628  
0 4632 4 1 2 4514 4579 
0 4633 4 1 2 4580 4511 
0 4634 4 2 2 4582 4583 
2 4635 1 4634  
2 4636 1 4634  
0 4637 4 3 2 4585 1204 
2 4638 1 4637  
2 4639 1 4637  
2 4640 1 4637  
0 4641 4 1 2 4523 4588 
0 4642 4 1 2 4589 1253 
0 4643 4 2 2 4404 4590 
2 4644 1 4643  
2 4645 1 4643  
0 4646 4 3 2 4593 4527 
2 4647 1 4646  
2 4648 1 4646  
2 4649 1 4646  
0 4650 4 3 2 4596 4532 
2 4651 1 4650  
2 4652 1 4650  
2 4653 1 4650  
0 4654 4 3 2 4599 4537 
2 4655 1 4654  
2 4656 1 4654  
2 4657 1 4654  
0 4658 4 3 2 4602 4542 
2 4659 1 4658  
2 4660 1 4658  
2 4661 1 4658  
0 4662 4 3 2 4605 4547 
2 4663 1 4662  
2 4664 1 4662  
2 4665 1 4662  
0 4666 4 1 2 4556 4608 
0 4667 4 1 2 4609 4553 
0 4668 4 2 2 4611 4612 
2 4669 1 4668  
2 4670 1 4668  
0 4671 4 3 2 4614 913 
2 4672 1 4671  
2 4673 1 4671  
2 4674 1 4671  
0 4675 4 1 2 4565 4617 
0 4676 4 1 2 4618 962 
0 4677 4 2 2 4438 4619 
2 4678 1 4677  
2 4679 1 4677  
0 4680 4 2 2 4620 4621 
2 4681 1 4680  
2 4682 1 4680  
0 4683 4 3 2 4626 4623 
2 4684 1 4683  
2 4685 1 4683  
2 4686 1 4683  
0 4687 4 1 2 4577 4629 
0 4688 4 1 2 4630 4574 
0 4689 4 2 2 4632 4633 
2 4690 1 4689  
2 4691 1 4689  
0 4692 4 3 2 4635 1156 
2 4693 1 4692  
2 4694 1 4692  
2 4695 1 4692  
0 4696 4 1 2 4586 4638 
0 4697 4 1 2 4639 1205 
0 4698 4 2 2 4459 4640 
2 4699 1 4698  
2 4700 1 4698  
0 4701 4 2 2 4641 4642 
2 4702 1 4701  
2 4703 1 4701  
0 4704 4 3 2 1300 4644 
2 4705 1 4704  
2 4706 1 4704  
2 4707 1 4704  
0 4708 4 1 2 4594 4647 
0 4709 4 1 2 4648 4528 
0 4710 4 1 2 4597 4651 
0 4711 4 1 2 4652 4533 
0 4712 4 1 2 4600 4655 
0 4713 4 1 2 4656 4538 
0 4714 4 1 2 4603 4659 
0 4715 4 1 2 4660 4543 
0 4716 4 1 2 4606 4663 
0 4717 4 1 2 4664 4548 
0 4718 4 2 2 4666 4667 
2 4719 1 4718  
2 4720 1 4718  
0 4721 4 3 2 4669 865 
2 4722 1 4721  
2 4723 1 4721  
2 4724 1 4721  
0 4725 4 1 2 4615 4672 
0 4726 4 1 2 4673 914 
0 4727 4 2 2 4497 4674 
2 4728 1 4727  
2 4729 1 4727  
0 4730 4 2 2 4675 4676 
2 4731 1 4730  
2 4732 1 4730  
0 4733 4 3 2 4681 4678 
2 4734 1 4733  
2 4735 1 4733  
2 4736 1 4733  
0 4737 4 1 2 4627 4684 
0 4738 4 1 2 4685 4624 
0 4739 4 2 2 4687 4688 
2 4740 1 4739  
2 4741 1 4739  
0 4742 4 3 2 4690 1108 
2 4743 1 4742  
2 4744 1 4742  
2 4745 1 4742  
0 4746 4 1 2 4636 4693 
0 4747 4 1 2 4694 1157 
0 4748 4 2 2 4518 4695 
2 4749 1 4748  
2 4750 1 4748  
0 4751 4 2 2 4696 4697 
2 4752 1 4751  
2 4753 1 4751  
0 4754 4 3 2 4702 4699 
2 4755 1 4754  
2 4756 1 4754  
2 4757 1 4754  
0 4758 4 1 2 1301 4705 
0 4759 4 1 2 4706 4645 
0 4760 4 2 2 4708 4709 
2 4761 1 4760  
2 4762 1 4760  
0 4763 4 2 2 4710 4711 
2 4764 1 4763  
2 4765 1 4763  
0 4766 4 2 2 4712 4713 
2 4767 1 4766  
2 4768 1 4766  
0 4769 4 2 2 4714 4715 
2 4770 1 4769  
2 4771 1 4769  
0 4772 4 2 2 4716 4717 
2 4773 1 4772  
2 4774 1 4772  
0 4775 4 3 2 4719 817 
2 4776 1 4775  
2 4777 1 4775  
2 4778 1 4775  
0 4779 4 1 2 4670 4722 
0 4780 4 1 2 4723 866 
0 4781 4 2 2 4560 4724 
2 4782 1 4781  
2 4783 1 4781  
0 4784 4 2 2 4725 4726 
2 4785 1 4784  
2 4786 1 4784  
0 4787 4 3 2 4731 4728 
2 4788 1 4787  
2 4789 1 4787  
2 4790 1 4787  
0 4791 4 1 2 4682 4734 
0 4792 4 1 2 4735 4679 
0 4793 4 2 2 4737 4738 
2 4794 1 4793  
2 4795 1 4793  
0 4796 4 3 2 4740 1060 
2 4797 1 4796  
2 4798 1 4796  
2 4799 1 4796  
0 4800 4 1 2 4691 4743 
0 4801 4 1 2 4744 1109 
0 4802 4 2 2 4581 4745 
2 4803 1 4802  
2 4804 1 4802  
0 4805 4 2 2 4746 4747 
2 4806 1 4805  
2 4807 1 4805  
0 4808 4 3 2 4752 4749 
2 4809 1 4808  
2 4810 1 4808  
2 4811 1 4808  
0 4812 4 1 2 4703 4755 
0 4813 4 1 2 4756 4700 
0 4814 4 2 2 4758 4759 
2 4815 1 4814  
2 4816 1 4814  
0 4817 4 3 2 4761 577 
2 4818 1 4817  
2 4819 1 4817  
2 4820 1 4817  
0 4821 4 3 2 4764 625 
2 4822 1 4821  
2 4823 1 4821  
2 4824 1 4821  
0 4825 4 3 2 4767 673 
2 4826 1 4825  
2 4827 1 4825  
2 4828 1 4825  
0 4829 4 3 2 4770 721 
2 4830 1 4829  
2 4831 1 4829  
2 4832 1 4829  
0 4833 4 3 2 4773 769 
2 4834 1 4833  
2 4835 1 4833  
2 4836 1 4833  
0 4837 4 1 2 4720 4776 
0 4838 4 1 2 4777 818 
0 4839 4 2 2 4610 4778 
2 4840 1 4839  
2 4841 1 4839  
0 4842 4 2 2 4779 4780 
2 4843 1 4842  
2 4844 1 4842  
0 4845 4 3 2 4785 4782 
2 4846 1 4845  
2 4847 1 4845  
2 4848 1 4845  
0 4849 4 1 2 4732 4788 
0 4850 4 1 2 4789 4729 
0 4851 4 2 2 4791 4792 
2 4852 1 4851  
2 4853 1 4851  
0 4854 4 3 2 4794 1012 
2 4855 1 4854  
2 4856 1 4854  
2 4857 1 4854  
0 4858 4 1 2 4741 4797 
0 4859 4 1 2 4798 1061 
0 4860 4 2 2 4631 4799 
2 4861 1 4860  
2 4862 1 4860  
0 4863 4 2 2 4800 4801 
2 4864 1 4863  
2 4865 1 4863  
0 4866 4 3 2 4806 4803 
2 4867 1 4866  
2 4868 1 4866  
2 4869 1 4866  
0 4870 4 1 2 4753 4809 
0 4871 4 1 2 4810 4750 
0 4872 4 2 2 4812 4813 
2 4873 1 4872  
2 4874 1 4872  
0 4875 4 3 2 4815 1255 
2 4876 1 4875  
2 4877 1 4875  
2 4878 1 4875  
0 4879 4 1 2 4762 4818 
0 4880 4 1 2 4819 578 
0 4881 4 2 2 4649 4820 
2 4882 1 4881  
2 4883 1 4881  
0 4884 4 1 2 4765 4822 
0 4885 4 1 2 4823 626 
0 4886 4 2 2 4653 4824 
2 4887 1 4886  
2 4888 1 4886  
0 4889 4 1 2 4768 4826 
0 4890 4 1 2 4827 674 
0 4891 4 2 2 4657 4828 
2 4892 1 4891  
2 4893 1 4891  
0 4894 4 1 2 4771 4830 
0 4895 4 1 2 4831 722 
0 4896 4 2 2 4661 4832 
2 4897 1 4896  
2 4898 1 4896  
0 4899 4 1 2 4774 4834 
0 4900 4 1 2 4835 770 
0 4901 4 2 2 4665 4836 
2 4902 1 4901  
2 4903 1 4901  
0 4904 4 2 2 4837 4838 
2 4905 1 4904  
2 4906 1 4904  
0 4907 4 3 2 4843 4840 
2 4908 1 4907  
2 4909 1 4907  
2 4910 1 4907  
0 4911 4 1 2 4786 4846 
0 4912 4 1 2 4847 4783 
0 4913 4 2 2 4849 4850 
2 4914 1 4913  
2 4915 1 4913  
0 4916 4 3 2 4852 964 
2 4917 1 4916  
2 4918 1 4916  
2 4919 1 4916  
0 4920 4 1 2 4795 4855 
0 4921 4 1 2 4856 1013 
0 4922 4 2 2 4686 4857 
2 4923 1 4922  
2 4924 1 4922  
0 4925 4 2 2 4858 4859 
2 4926 1 4925  
2 4927 1 4925  
0 4928 4 3 2 4864 4861 
2 4929 1 4928  
2 4930 1 4928  
2 4931 1 4928  
0 4932 4 1 2 4807 4867 
0 4933 4 1 2 4868 4804 
0 4934 4 2 2 4870 4871 
2 4935 1 4934  
2 4936 1 4934  
0 4937 4 3 2 4873 1207 
2 4938 1 4937  
2 4939 1 4937  
2 4940 1 4937  
0 4941 4 1 2 4816 4876 
0 4942 4 1 2 4877 1256 
0 4943 4 2 2 4707 4878 
2 4944 1 4943  
2 4945 1 4943  
3 4946 4 0 2 4879 4880 
0 4947 4 2 2 4884 4885 
2 4948 1 4947  
2 4949 1 4947  
0 4950 4 2 2 4889 4890 
2 4951 1 4950  
2 4952 1 4950  
0 4953 4 2 2 4894 4895 
2 4954 1 4953  
2 4955 1 4953  
0 4956 4 2 2 4899 4900 
2 4957 1 4956  
2 4958 1 4956  
0 4959 4 3 2 4905 4902 
2 4960 1 4959  
2 4961 1 4959  
2 4962 1 4959  
0 4963 4 1 2 4844 4908 
0 4964 4 1 2 4909 4841 
0 4965 4 2 2 4911 4912 
2 4966 1 4965  
2 4967 1 4965  
0 4968 4 3 2 4914 916 
2 4969 1 4968  
2 4970 1 4968  
2 4971 1 4968  
0 4972 4 1 2 4853 4917 
0 4973 4 1 2 4918 965 
0 4974 4 2 2 4736 4919 
2 4975 1 4974  
2 4976 1 4974  
0 4977 4 2 2 4920 4921 
2 4978 1 4977  
2 4979 1 4977  
0 4980 4 3 2 4926 4923 
2 4981 1 4980  
2 4982 1 4980  
2 4983 1 4980  
0 4984 4 1 2 4865 4929 
0 4985 4 1 2 4930 4862 
0 4986 4 2 2 4932 4933 
2 4987 1 4986  
2 4988 1 4986  
0 4989 4 3 2 4935 1159 
2 4990 1 4989  
2 4991 1 4989  
2 4992 1 4989  
0 4993 4 1 2 4874 4938 
0 4994 4 1 2 4939 1208 
0 4995 4 2 2 4757 4940 
2 4996 1 4995  
2 4997 1 4995  
0 4998 4 2 2 4941 4942 
2 4999 1 4998  
2 5000 1 4998  
0 5001 4 3 2 1303 4944 
2 5002 1 5001  
2 5003 1 5001  
2 5004 1 5001  
0 5005 4 3 2 4948 4882 
2 5006 1 5005  
2 5007 1 5005  
2 5008 1 5005  
0 5009 4 3 2 4951 4887 
2 5010 1 5009  
2 5011 1 5009  
2 5012 1 5009  
0 5013 4 3 2 4954 4892 
2 5014 1 5013  
2 5015 1 5013  
2 5016 1 5013  
0 5017 4 3 2 4957 4897 
2 5018 1 5017  
2 5019 1 5017  
2 5020 1 5017  
0 5021 4 1 2 4906 4960 
0 5022 4 1 2 4961 4903 
0 5023 4 2 2 4963 4964 
2 5024 1 5023  
2 5025 1 5023  
0 5026 4 3 2 4966 868 
2 5027 1 5026  
2 5028 1 5026  
2 5029 1 5026  
0 5030 4 1 2 4915 4969 
0 5031 4 1 2 4970 917 
0 5032 4 2 2 4790 4971 
2 5033 1 5032  
2 5034 1 5032  
0 5035 4 2 2 4972 4973 
2 5036 1 5035  
2 5037 1 5035  
0 5038 4 3 2 4978 4975 
2 5039 1 5038  
2 5040 1 5038  
2 5041 1 5038  
0 5042 4 1 2 4927 4981 
0 5043 4 1 2 4982 4924 
0 5044 4 2 2 4984 4985 
2 5045 1 5044  
2 5046 1 5044  
0 5047 4 3 2 4987 1111 
2 5048 1 5047  
2 5049 1 5047  
2 5050 1 5047  
0 5051 4 1 2 4936 4990 
0 5052 4 1 2 4991 1160 
0 5053 4 2 2 4811 4992 
2 5054 1 5053  
2 5055 1 5053  
0 5056 4 2 2 4993 4994 
2 5057 1 5056  
2 5058 1 5056  
0 5059 4 3 2 4999 4996 
2 5060 1 5059  
2 5061 1 5059  
2 5062 1 5059  
0 5063 4 1 2 1304 5002 
0 5064 4 1 2 5003 4945 
0 5065 4 1 2 4949 5006 
0 5066 4 1 2 5007 4883 
0 5067 4 1 2 4952 5010 
0 5068 4 1 2 5011 4888 
0 5069 4 1 2 4955 5014 
0 5070 4 1 2 5015 4893 
0 5071 4 1 2 4958 5018 
0 5072 4 1 2 5019 4898 
0 5073 4 2 2 5021 5022 
2 5074 1 5073  
2 5075 1 5073  
0 5076 4 3 2 5024 820 
2 5077 1 5076  
2 5078 1 5076  
2 5079 1 5076  
0 5080 4 1 2 4967 5027 
0 5081 4 1 2 5028 869 
0 5082 4 2 2 4848 5029 
2 5083 1 5082  
2 5084 1 5082  
0 5085 4 2 2 5030 5031 
2 5086 1 5085  
2 5087 1 5085  
0 5088 4 3 2 5036 5033 
2 5089 1 5088  
2 5090 1 5088  
2 5091 1 5088  
0 5092 4 1 2 4979 5039 
0 5093 4 1 2 5040 4976 
0 5094 4 2 2 5042 5043 
2 5095 1 5094  
2 5096 1 5094  
0 5097 4 3 2 5045 1063 
2 5098 1 5097  
2 5099 1 5097  
2 5100 1 5097  
0 5101 4 1 2 4988 5048 
0 5102 4 1 2 5049 1112 
0 5103 4 2 2 4869 5050 
2 5104 1 5103  
2 5105 1 5103  
0 5106 4 2 2 5051 5052 
2 5107 1 5106  
2 5108 1 5106  
0 5109 4 3 2 5057 5054 
2 5110 1 5109  
2 5111 1 5109  
2 5112 1 5109  
0 5113 4 1 2 5000 5060 
0 5114 4 1 2 5061 4997 
0 5115 4 2 2 5063 5064 
2 5116 1 5115  
2 5117 1 5115  
0 5118 4 2 2 5065 5066 
2 5119 1 5118  
2 5120 1 5118  
0 5121 4 2 2 5067 5068 
2 5122 1 5121  
2 5123 1 5121  
0 5124 4 2 2 5069 5070 
2 5125 1 5124  
2 5126 1 5124  
0 5127 4 2 2 5071 5072 
2 5128 1 5127  
2 5129 1 5127  
0 5130 4 3 2 5074 772 
2 5131 1 5130  
2 5132 1 5130  
2 5133 1 5130  
0 5134 4 1 2 5025 5077 
0 5135 4 1 2 5078 821 
0 5136 4 2 2 4910 5079 
2 5137 1 5136  
2 5138 1 5136  
0 5139 4 2 2 5080 5081 
2 5140 1 5139  
2 5141 1 5139  
0 5142 4 3 2 5086 5083 
2 5143 1 5142  
2 5144 1 5142  
2 5145 1 5142  
0 5146 4 1 2 5037 5089 
0 5147 4 1 2 5090 5034 
0 5148 4 2 2 5092 5093 
2 5149 1 5148  
2 5150 1 5148  
0 5151 4 3 2 5095 1015 
2 5152 1 5151  
2 5153 1 5151  
2 5154 1 5151  
0 5155 4 1 2 5046 5098 
0 5156 4 1 2 5099 1064 
0 5157 4 2 2 4931 5100 
2 5158 1 5157  
2 5159 1 5157  
0 5160 4 2 2 5101 5102 
2 5161 1 5160  
2 5162 1 5160  
0 5163 4 3 2 5107 5104 
2 5164 1 5163  
2 5165 1 5163  
2 5166 1 5163  
0 5167 4 1 2 5058 5110 
0 5168 4 1 2 5111 5055 
0 5169 4 2 2 5113 5114 
2 5170 1 5169  
2 5171 1 5169  
0 5172 4 3 2 5116 1258 
2 5173 1 5172  
2 5174 1 5172  
2 5175 1 5172  
0 5176 4 3 2 5119 580 
2 5177 1 5176  
2 5178 1 5176  
2 5179 1 5176  
0 5180 4 3 2 5122 628 
2 5181 1 5180  
2 5182 1 5180  
2 5183 1 5180  
0 5184 4 3 2 5125 676 
2 5185 1 5184  
2 5186 1 5184  
2 5187 1 5184  
0 5188 4 3 2 5128 724 
2 5189 1 5188  
2 5190 1 5188  
2 5191 1 5188  
0 5192 4 1 2 5075 5131 
0 5193 4 1 2 5132 773 
0 5194 4 2 2 4962 5133 
2 5195 1 5194  
2 5196 1 5194  
0 5197 4 2 2 5134 5135 
2 5198 1 5197  
2 5199 1 5197  
0 5200 4 3 2 5140 5137 
2 5201 1 5200  
2 5202 1 5200  
2 5203 1 5200  
0 5204 4 1 2 5087 5143 
0 5205 4 1 2 5144 5084 
0 5206 4 2 2 5146 5147 
2 5207 1 5206  
2 5208 1 5206  
0 5209 4 3 2 5149 967 
2 5210 1 5209  
2 5211 1 5209  
2 5212 1 5209  
0 5213 4 1 2 5096 5152 
0 5214 4 1 2 5153 1016 
0 5215 4 2 2 4983 5154 
2 5216 1 5215  
2 5217 1 5215  
0 5218 4 2 2 5155 5156 
2 5219 1 5218  
2 5220 1 5218  
0 5221 4 3 2 5161 5158 
2 5222 1 5221  
2 5223 1 5221  
2 5224 1 5221  
0 5225 4 1 2 5108 5164 
0 5226 4 1 2 5165 5105 
0 5227 4 2 2 5167 5168 
2 5228 1 5227  
2 5229 1 5227  
0 5230 4 3 2 5170 1210 
2 5231 1 5230  
2 5232 1 5230  
2 5233 1 5230  
0 5234 4 1 2 5117 5173 
0 5235 4 1 2 5174 1259 
0 5236 4 2 2 5004 5175 
2 5237 1 5236  
2 5238 1 5236  
0 5239 4 1 2 5120 5177 
0 5240 4 1 2 5178 581 
0 5241 4 2 2 5008 5179 
2 5242 1 5241  
2 5243 1 5241  
0 5244 4 1 2 5123 5181 
0 5245 4 1 2 5182 629 
0 5246 4 2 2 5012 5183 
2 5247 1 5246  
2 5248 1 5246  
0 5249 4 1 2 5126 5185 
0 5250 4 1 2 5186 677 
0 5251 4 2 2 5016 5187 
2 5252 1 5251  
2 5253 1 5251  
0 5254 4 1 2 5129 5189 
0 5255 4 1 2 5190 725 
0 5256 4 2 2 5020 5191 
2 5257 1 5256  
2 5258 1 5256  
0 5259 4 2 2 5192 5193 
2 5260 1 5259  
2 5261 1 5259  
0 5262 4 3 2 5198 5195 
2 5263 1 5262  
2 5264 1 5262  
2 5265 1 5262  
0 5266 4 1 2 5141 5201 
0 5267 4 1 2 5202 5138 
0 5268 4 2 2 5204 5205 
2 5269 1 5268  
2 5270 1 5268  
0 5271 4 3 2 5207 919 
2 5272 1 5271  
2 5273 1 5271  
2 5274 1 5271  
0 5275 4 1 2 5150 5210 
0 5276 4 1 2 5211 968 
0 5277 4 2 2 5041 5212 
2 5278 1 5277  
2 5279 1 5277  
0 5280 4 2 2 5213 5214 
2 5281 1 5280  
2 5282 1 5280  
0 5283 4 3 2 5219 5216 
2 5284 1 5283  
2 5285 1 5283  
2 5286 1 5283  
0 5287 4 1 2 5162 5222 
0 5288 4 1 2 5223 5159 
0 5289 4 2 2 5225 5226 
2 5290 1 5289  
2 5291 1 5289  
0 5292 4 3 2 5228 1162 
2 5293 1 5292  
2 5294 1 5292  
2 5295 1 5292  
0 5296 4 1 2 5171 5231 
0 5297 4 1 2 5232 1211 
0 5298 4 2 2 5062 5233 
2 5299 1 5298  
2 5300 1 5298  
0 5301 4 2 2 5234 5235 
2 5302 1 5301  
2 5303 1 5301  
0 5304 4 3 2 1306 5237 
2 5305 1 5304  
2 5306 1 5304  
2 5307 1 5304  
3 5308 4 0 2 5239 5240 
0 5309 4 2 2 5244 5245 
2 5310 1 5309  
2 5311 1 5309  
0 5312 4 2 2 5249 5250 
2 5313 1 5312  
2 5314 1 5312  
0 5315 4 2 2 5254 5255 
2 5316 1 5315  
2 5317 1 5315  
0 5318 4 3 2 5260 5257 
2 5319 1 5318  
2 5320 1 5318  
2 5321 1 5318  
0 5322 4 1 2 5199 5263 
0 5323 4 1 2 5264 5196 
0 5324 4 2 2 5266 5267 
2 5325 1 5324  
2 5326 1 5324  
0 5327 4 3 2 5269 871 
2 5328 1 5327  
2 5329 1 5327  
2 5330 1 5327  
0 5331 4 1 2 5208 5272 
0 5332 4 1 2 5273 920 
0 5333 4 2 2 5091 5274 
2 5334 1 5333  
2 5335 1 5333  
0 5336 4 2 2 5275 5276 
2 5337 1 5336  
2 5338 1 5336  
0 5339 4 3 2 5281 5278 
2 5340 1 5339  
2 5341 1 5339  
2 5342 1 5339  
0 5343 4 1 2 5220 5284 
0 5344 4 1 2 5285 5217 
0 5345 4 2 2 5287 5288 
2 5346 1 5345  
2 5347 1 5345  
0 5348 4 3 2 5290 1114 
2 5349 1 5348  
2 5350 1 5348  
2 5351 1 5348  
0 5352 4 1 2 5229 5293 
0 5353 4 1 2 5294 1163 
0 5354 4 2 2 5112 5295 
2 5355 1 5354  
2 5356 1 5354  
0 5357 4 2 2 5296 5297 
2 5358 1 5357  
2 5359 1 5357  
0 5360 4 3 2 5302 5299 
2 5361 1 5360  
2 5362 1 5360  
2 5363 1 5360  
0 5364 4 1 2 1307 5305 
0 5365 4 1 2 5306 5238 
0 5366 4 3 2 5310 5242 
2 5367 1 5366  
2 5368 1 5366  
2 5369 1 5366  
0 5370 4 3 2 5313 5247 
2 5371 1 5370  
2 5372 1 5370  
2 5373 1 5370  
0 5374 4 3 2 5316 5252 
2 5375 1 5374  
2 5376 1 5374  
2 5377 1 5374  
0 5378 4 1 2 5261 5319 
0 5379 4 1 2 5320 5258 
0 5380 4 2 2 5322 5323 
2 5381 1 5380  
2 5382 1 5380  
0 5383 4 3 2 5325 823 
2 5384 1 5383  
2 5385 1 5383  
2 5386 1 5383  
0 5387 4 1 2 5270 5328 
0 5388 4 1 2 5329 872 
0 5389 4 2 2 5145 5330 
2 5390 1 5389  
2 5391 1 5389  
0 5392 4 2 2 5331 5332 
2 5393 1 5392  
2 5394 1 5392  
0 5395 4 3 2 5337 5334 
2 5396 1 5395  
2 5397 1 5395  
2 5398 1 5395  
0 5399 4 1 2 5282 5340 
0 5400 4 1 2 5341 5279 
0 5401 4 2 2 5343 5344 
2 5402 1 5401  
2 5403 1 5401  
0 5404 4 3 2 5346 1066 
2 5405 1 5404  
2 5406 1 5404  
2 5407 1 5404  
0 5408 4 1 2 5291 5349 
0 5409 4 1 2 5350 1115 
0 5410 4 2 2 5166 5351 
2 5411 1 5410  
2 5412 1 5410  
0 5413 4 2 2 5352 5353 
2 5414 1 5413  
2 5415 1 5413  
0 5416 4 3 2 5358 5355 
2 5417 1 5416  
2 5418 1 5416  
2 5419 1 5416  
0 5420 4 1 2 5303 5361 
0 5421 4 1 2 5362 5300 
0 5422 4 2 2 5364 5365 
2 5423 1 5422  
2 5424 1 5422  
0 5425 4 1 2 5311 5367 
0 5426 4 1 2 5368 5243 
0 5427 4 1 2 5314 5371 
0 5428 4 1 2 5372 5248 
0 5429 4 1 2 5317 5375 
0 5430 4 1 2 5376 5253 
0 5431 4 2 2 5378 5379 
2 5432 1 5431  
2 5433 1 5431  
0 5434 4 3 2 5381 775 
2 5435 1 5434  
2 5436 1 5434  
2 5437 1 5434  
0 5438 4 1 2 5326 5384 
0 5439 4 1 2 5385 824 
0 5440 4 2 2 5203 5386 
2 5441 1 5440  
2 5442 1 5440  
0 5443 4 2 2 5387 5388 
2 5444 1 5443  
2 5445 1 5443  
0 5446 4 3 2 5393 5390 
2 5447 1 5446  
2 5448 1 5446  
2 5449 1 5446  
0 5450 4 1 2 5338 5396 
0 5451 4 1 2 5397 5335 
0 5452 4 2 2 5399 5400 
2 5453 1 5452  
2 5454 1 5452  
0 5455 4 3 2 5402 1018 
2 5456 1 5455  
2 5457 1 5455  
2 5458 1 5455  
0 5459 4 1 2 5347 5405 
0 5460 4 1 2 5406 1067 
0 5461 4 2 2 5224 5407 
2 5462 1 5461  
2 5463 1 5461  
0 5464 4 2 2 5408 5409 
2 5465 1 5464  
2 5466 1 5464  
0 5467 4 3 2 5414 5411 
2 5468 1 5467  
2 5469 1 5467  
2 5470 1 5467  
0 5471 4 1 2 5359 5417 
0 5472 4 1 2 5418 5356 
0 5473 4 2 2 5420 5421 
2 5474 1 5473  
2 5475 1 5473  
0 5476 4 3 2 5423 1261 
2 5477 1 5476  
2 5478 1 5476  
2 5479 1 5476  
0 5480 4 2 2 5425 5426 
2 5481 1 5480  
2 5482 1 5480  
0 5483 4 2 2 5427 5428 
2 5484 1 5483  
2 5485 1 5483  
0 5486 4 2 2 5429 5430 
2 5487 1 5486  
2 5488 1 5486  
0 5489 4 3 2 5432 727 
2 5490 1 5489  
2 5491 1 5489  
2 5492 1 5489  
0 5493 4 1 2 5382 5435 
0 5494 4 1 2 5436 776 
0 5495 4 2 2 5265 5437 
2 5496 1 5495  
2 5497 1 5495  
0 5498 4 2 2 5438 5439 
2 5499 1 5498  
2 5500 1 5498  
0 5501 4 3 2 5444 5441 
2 5502 1 5501  
2 5503 1 5501  
2 5504 1 5501  
0 5505 4 1 2 5394 5447 
0 5506 4 1 2 5448 5391 
0 5507 4 2 2 5450 5451 
2 5508 1 5507  
2 5509 1 5507  
0 5510 4 3 2 5453 970 
2 5511 1 5510  
2 5512 1 5510  
2 5513 1 5510  
0 5514 4 1 2 5403 5456 
0 5515 4 1 2 5457 1019 
0 5516 4 2 2 5286 5458 
2 5517 1 5516  
2 5518 1 5516  
0 5519 4 2 2 5459 5460 
2 5520 1 5519  
2 5521 1 5519  
0 5522 4 3 2 5465 5462 
2 5523 1 5522  
2 5524 1 5522  
2 5525 1 5522  
0 5526 4 1 2 5415 5468 
0 5527 4 1 2 5469 5412 
0 5528 4 2 2 5471 5472 
2 5529 1 5528  
2 5530 1 5528  
0 5531 4 3 2 5474 1213 
2 5532 1 5531  
2 5533 1 5531  
2 5534 1 5531  
0 5535 4 1 2 5424 5477 
0 5536 4 1 2 5478 1262 
0 5537 4 2 2 5307 5479 
2 5538 1 5537  
2 5539 1 5537  
0 5540 4 3 2 5481 583 
2 5541 1 5540  
2 5542 1 5540  
2 5543 1 5540  
0 5544 4 3 2 5484 631 
2 5545 1 5544  
2 5546 1 5544  
2 5547 1 5544  
0 5548 4 3 2 5487 679 
2 5549 1 5548  
2 5550 1 5548  
2 5551 1 5548  
0 5552 4 1 2 5433 5490 
0 5553 4 1 2 5491 728 
0 5554 4 2 2 5321 5492 
2 5555 1 5554  
2 5556 1 5554  
0 5557 4 2 2 5493 5494 
2 5558 1 5557  
2 5559 1 5557  
0 5560 4 3 2 5499 5496 
2 5561 1 5560  
2 5562 1 5560  
2 5563 1 5560  
0 5564 4 1 2 5445 5502 
0 5565 4 1 2 5503 5442 
0 5566 4 2 2 5505 5506 
2 5567 1 5566  
2 5568 1 5566  
0 5569 4 3 2 5508 922 
2 5570 1 5569  
2 5571 1 5569  
2 5572 1 5569  
0 5573 4 1 2 5454 5511 
0 5574 4 1 2 5512 971 
0 5575 4 2 2 5342 5513 
2 5576 1 5575  
2 5577 1 5575  
0 5578 4 2 2 5514 5515 
2 5579 1 5578  
2 5580 1 5578  
0 5581 4 3 2 5520 5517 
2 5582 1 5581  
2 5583 1 5581  
2 5584 1 5581  
0 5585 4 1 2 5466 5523 
0 5586 4 1 2 5524 5463 
0 5587 4 2 2 5526 5527 
2 5588 1 5587  
2 5589 1 5587  
0 5590 4 3 2 5529 1165 
2 5591 1 5590  
2 5592 1 5590  
2 5593 1 5590  
0 5594 4 1 2 5475 5532 
0 5595 4 1 2 5533 1214 
0 5596 4 2 2 5363 5534 
2 5597 1 5596  
2 5598 1 5596  
0 5599 4 2 2 5535 5536 
2 5600 1 5599  
2 5601 1 5599  
0 5602 4 3 2 1309 5538 
2 5603 1 5602  
2 5604 1 5602  
2 5605 1 5602  
0 5606 4 1 2 5482 5541 
0 5607 4 1 2 5542 584 
0 5608 4 2 2 5369 5543 
2 5609 1 5608  
2 5610 1 5608  
0 5611 4 1 2 5485 5545 
0 5612 4 1 2 5546 632 
0 5613 4 2 2 5373 5547 
2 5614 1 5613  
2 5615 1 5613  
0 5616 4 1 2 5488 5549 
0 5617 4 1 2 5550 680 
0 5618 4 2 2 5377 5551 
2 5619 1 5618  
2 5620 1 5618  
0 5621 4 2 2 5552 5553 
2 5622 1 5621  
2 5623 1 5621  
0 5624 4 3 2 5558 5555 
2 5625 1 5624  
2 5626 1 5624  
2 5627 1 5624  
0 5628 4 1 2 5500 5561 
0 5629 4 1 2 5562 5497 
0 5630 4 2 2 5564 5565 
2 5631 1 5630  
2 5632 1 5630  
0 5633 4 3 2 5567 874 
2 5634 1 5633  
2 5635 1 5633  
2 5636 1 5633  
0 5637 4 1 2 5509 5570 
0 5638 4 1 2 5571 923 
0 5639 4 2 2 5398 5572 
2 5640 1 5639  
2 5641 1 5639  
0 5642 4 2 2 5573 5574 
2 5643 1 5642  
2 5644 1 5642  
0 5645 4 3 2 5579 5576 
2 5646 1 5645  
2 5647 1 5645  
2 5648 1 5645  
0 5649 4 1 2 5521 5582 
0 5650 4 1 2 5583 5518 
0 5651 4 2 2 5585 5586 
2 5652 1 5651  
2 5653 1 5651  
0 5654 4 3 2 5588 1117 
2 5655 1 5654  
2 5656 1 5654  
2 5657 1 5654  
0 5658 4 1 2 5530 5591 
0 5659 4 1 2 5592 1166 
0 5660 4 2 2 5419 5593 
2 5661 1 5660  
2 5662 1 5660  
0 5663 4 2 2 5594 5595 
2 5664 1 5663  
2 5665 1 5663  
0 5666 4 3 2 5600 5597 
2 5667 1 5666  
2 5668 1 5666  
2 5669 1 5666  
0 5670 4 1 2 1310 5603 
0 5671 4 1 2 5604 5539 
3 5672 4 0 2 5606 5607 
0 5673 4 2 2 5611 5612 
2 5674 1 5673  
2 5675 1 5673  
0 5676 4 2 2 5616 5617 
2 5677 1 5676  
2 5678 1 5676  
0 5679 4 3 2 5622 5619 
2 5680 1 5679  
2 5681 1 5679  
2 5682 1 5679  
0 5683 4 1 2 5559 5625 
0 5684 4 1 2 5626 5556 
0 5685 4 2 2 5628 5629 
2 5686 1 5685  
2 5687 1 5685  
0 5688 4 3 2 5631 826 
2 5689 1 5688  
2 5690 1 5688  
2 5691 1 5688  
0 5692 4 1 2 5568 5634 
0 5693 4 1 2 5635 875 
0 5694 4 2 2 5449 5636 
2 5695 1 5694  
2 5696 1 5694  
0 5697 4 2 2 5637 5638 
2 5698 1 5697  
2 5699 1 5697  
0 5700 4 3 2 5643 5640 
2 5701 1 5700  
2 5702 1 5700  
2 5703 1 5700  
0 5704 4 1 2 5580 5646 
0 5705 4 1 2 5647 5577 
0 5706 4 2 2 5649 5650 
2 5707 1 5706  
2 5708 1 5706  
0 5709 4 3 2 5652 1069 
2 5710 1 5709  
2 5711 1 5709  
2 5712 1 5709  
0 5713 4 1 2 5589 5655 
0 5714 4 1 2 5656 1118 
0 5715 4 2 2 5470 5657 
2 5716 1 5715  
2 5717 1 5715  
0 5718 4 2 2 5658 5659 
2 5719 1 5718  
2 5720 1 5718  
0 5721 4 3 2 5664 5661 
2 5722 1 5721  
2 5723 1 5721  
2 5724 1 5721  
0 5725 4 1 2 5601 5667 
0 5726 4 1 2 5668 5598 
0 5727 4 2 2 5670 5671 
2 5728 1 5727  
2 5729 1 5727  
0 5730 4 3 2 5674 5609 
2 5731 1 5730  
2 5732 1 5730  
2 5733 1 5730  
0 5734 4 3 2 5677 5614 
2 5735 1 5734  
2 5736 1 5734  
2 5737 1 5734  
0 5738 4 1 2 5623 5680 
0 5739 4 1 2 5681 5620 
0 5740 4 2 2 5683 5684 
2 5741 1 5740  
2 5742 1 5740  
0 5743 4 3 2 5686 778 
2 5744 1 5743  
2 5745 1 5743  
2 5746 1 5743  
0 5747 4 1 2 5632 5689 
0 5748 4 1 2 5690 827 
0 5749 4 2 2 5504 5691 
2 5750 1 5749  
2 5751 1 5749  
0 5752 4 2 2 5692 5693 
2 5753 1 5752  
2 5754 1 5752  
0 5755 4 3 2 5698 5695 
2 5756 1 5755  
2 5757 1 5755  
2 5758 1 5755  
0 5759 4 1 2 5644 5701 
0 5760 4 1 2 5702 5641 
0 5761 4 2 2 5704 5705 
2 5762 1 5761  
2 5763 1 5761  
0 5764 4 3 2 5707 1021 
2 5765 1 5764  
2 5766 1 5764  
2 5767 1 5764  
0 5768 4 1 2 5653 5710 
0 5769 4 1 2 5711 1070 
0 5770 4 2 2 5525 5712 
2 5771 1 5770  
2 5772 1 5770  
0 5773 4 2 2 5713 5714 
2 5774 1 5773  
2 5775 1 5773  
0 5776 4 3 2 5719 5716 
2 5777 1 5776  
2 5778 1 5776  
2 5779 1 5776  
0 5780 4 1 2 5665 5722 
0 5781 4 1 2 5723 5662 
0 5782 4 2 2 5725 5726 
2 5783 1 5782  
2 5784 1 5782  
0 5785 4 1 2 5675 5731 
0 5786 4 1 2 5732 5610 
0 5787 4 1 2 5678 5735 
0 5788 4 1 2 5736 5615 
0 5789 4 2 2 5738 5739 
2 5790 1 5789  
2 5791 1 5789  
0 5792 4 3 2 5741 730 
2 5793 1 5792  
2 5794 1 5792  
2 5795 1 5792  
0 5796 4 1 2 5687 5744 
0 5797 4 1 2 5745 779 
0 5798 4 2 2 5563 5746 
2 5799 1 5798  
2 5800 1 5798  
0 5801 4 2 2 5747 5748 
2 5802 1 5801  
2 5803 1 5801  
0 5804 4 3 2 5753 5750 
2 5805 1 5804  
2 5806 1 5804  
2 5807 1 5804  
0 5808 4 1 2 5699 5756 
0 5809 4 1 2 5757 5696 
0 5810 4 2 2 5759 5760 
2 5811 1 5810  
2 5812 1 5810  
0 5813 4 3 2 5762 973 
2 5814 1 5813  
2 5815 1 5813  
2 5816 1 5813  
0 5817 4 1 2 5708 5765 
0 5818 4 1 2 5766 1022 
0 5819 4 2 2 5584 5767 
2 5820 1 5819  
2 5821 1 5819  
0 5822 4 2 2 5768 5769 
2 5823 1 5822  
2 5824 1 5822  
0 5825 4 3 2 5774 5771 
2 5826 1 5825  
2 5827 1 5825  
2 5828 1 5825  
0 5829 4 1 2 5720 5777 
0 5830 4 1 2 5778 5717 
0 5831 4 2 2 5780 5781 
2 5832 1 5831  
2 5833 1 5831  
0 5834 4 2 2 5785 5786 
2 5835 1 5834  
2 5836 1 5834  
0 5837 4 2 2 5787 5788 
2 5838 1 5837  
2 5839 1 5837  
0 5840 4 3 2 5790 682 
2 5841 1 5840  
2 5842 1 5840  
2 5843 1 5840  
0 5844 4 1 2 5742 5793 
0 5845 4 1 2 5794 731 
0 5846 4 2 2 5627 5795 
2 5847 1 5846  
2 5848 1 5846  
0 5849 4 2 2 5796 5797 
2 5850 1 5849  
2 5851 1 5849  
0 5852 4 3 2 5802 5799 
2 5853 1 5852  
2 5854 1 5852  
2 5855 1 5852  
0 5856 4 1 2 5754 5805 
0 5857 4 1 2 5806 5751 
0 5858 4 2 2 5808 5809 
2 5859 1 5858  
2 5860 1 5858  
0 5861 4 3 2 5811 925 
2 5862 1 5861  
2 5863 1 5861  
2 5864 1 5861  
0 5865 4 1 2 5763 5814 
0 5866 4 1 2 5815 974 
0 5867 4 2 2 5648 5816 
2 5868 1 5867  
2 5869 1 5867  
0 5870 4 2 2 5817 5818 
2 5871 1 5870  
2 5872 1 5870  
0 5873 4 3 2 5823 5820 
2 5874 1 5873  
2 5875 1 5873  
2 5876 1 5873  
0 5877 4 1 2 5775 5826 
0 5878 4 1 2 5827 5772 
0 5879 4 2 2 5829 5830 
2 5880 1 5879  
2 5881 1 5879  
0 5882 4 3 2 5835 586 
2 5883 1 5882  
2 5884 1 5882  
2 5885 1 5882  
0 5886 4 3 2 5838 634 
2 5887 1 5886  
2 5888 1 5886  
2 5889 1 5886  
0 5890 4 1 2 5791 5841 
0 5891 4 1 2 5842 683 
0 5892 4 2 2 5682 5843 
2 5893 1 5892  
2 5894 1 5892  
0 5895 4 2 2 5844 5845 
2 5896 1 5895  
2 5897 1 5895  
0 5898 4 3 2 5850 5847 
2 5899 1 5898  
2 5900 1 5898  
2 5901 1 5898  
0 5902 4 1 2 5803 5853 
0 5903 4 1 2 5854 5800 
0 5904 4 2 2 5856 5857 
2 5905 1 5904  
2 5906 1 5904  
0 5907 4 3 2 5859 877 
2 5908 1 5907  
2 5909 1 5907  
2 5910 1 5907  
0 5911 4 1 2 5812 5862 
0 5912 4 1 2 5863 926 
0 5913 4 2 2 5703 5864 
2 5914 1 5913  
2 5915 1 5913  
0 5916 4 2 2 5865 5866 
2 5917 1 5916  
2 5918 1 5916  
0 5919 4 3 2 5871 5868 
2 5920 1 5919  
2 5921 1 5919  
2 5922 1 5919  
0 5923 4 1 2 5824 5874 
0 5924 4 1 2 5875 5821 
0 5925 4 2 2 5877 5878 
2 5926 1 5925  
2 5927 1 5925  
0 5928 4 1 2 5836 5883 
0 5929 4 1 2 5884 587 
0 5930 4 2 2 5733 5885 
2 5931 1 5930  
2 5932 1 5930  
0 5933 4 1 2 5839 5887 
0 5934 4 1 2 5888 635 
0 5935 4 2 2 5737 5889 
2 5936 1 5935  
2 5937 1 5935  
0 5938 4 2 2 5890 5891 
2 5939 1 5938  
2 5940 1 5938  
0 5941 4 3 2 5896 5893 
2 5942 1 5941  
2 5943 1 5941  
2 5944 1 5941  
0 5945 4 1 2 5851 5899 
0 5946 4 1 2 5900 5848 
0 5947 4 2 2 5902 5903 
2 5948 1 5947  
2 5949 1 5947  
0 5950 4 3 2 5905 829 
2 5951 1 5950  
2 5952 1 5950  
2 5953 1 5950  
0 5954 4 1 2 5860 5908 
0 5955 4 1 2 5909 878 
0 5956 4 2 2 5758 5910 
2 5957 1 5956  
2 5958 1 5956  
0 5959 4 2 2 5911 5912 
2 5960 1 5959  
2 5961 1 5959  
0 5962 4 3 2 5917 5914 
2 5963 1 5962  
2 5964 1 5962  
2 5965 1 5962  
0 5966 4 1 2 5872 5920 
0 5967 4 1 2 5921 5869 
0 5968 4 2 2 5923 5924 
2 5969 1 5968  
2 5970 1 5968  
3 5971 4 0 2 5928 5929 
0 5972 4 2 2 5933 5934 
2 5973 1 5972  
2 5974 1 5972  
0 5975 4 3 2 5939 5936 
2 5976 1 5975  
2 5977 1 5975  
2 5978 1 5975  
0 5979 4 1 2 5897 5942 
0 5980 4 1 2 5943 5894 
0 5981 4 2 2 5945 5946 
2 5982 1 5981  
2 5983 1 5981  
0 5984 4 3 2 5948 781 
2 5985 1 5984  
2 5986 1 5984  
2 5987 1 5984  
0 5988 4 1 2 5906 5951 
0 5989 4 1 2 5952 830 
0 5990 4 2 2 5807 5953 
2 5991 1 5990  
2 5992 1 5990  
0 5993 4 2 2 5954 5955 
2 5994 1 5993  
2 5995 1 5993  
0 5996 4 3 2 5960 5957 
2 5997 1 5996  
2 5998 1 5996  
2 5999 1 5996  
0 6000 4 1 2 5918 5963 
0 6001 4 1 2 5964 5915 
0 6002 4 2 2 5966 5967 
2 6003 1 6002  
2 6004 1 6002  
0 6005 4 3 2 5973 5931 
2 6006 1 6005  
2 6007 1 6005  
2 6008 1 6005  
0 6009 4 1 2 5940 5976 
0 6010 4 1 2 5977 5937 
0 6011 4 2 2 5979 5980 
2 6012 1 6011  
2 6013 1 6011  
0 6014 4 3 2 5982 733 
2 6015 1 6014  
2 6016 1 6014  
2 6017 1 6014  
0 6018 4 1 2 5949 5985 
0 6019 4 1 2 5986 782 
0 6020 4 2 2 5855 5987 
2 6021 1 6020  
2 6022 1 6020  
0 6023 4 2 2 5988 5989 
2 6024 1 6023  
2 6025 1 6023  
0 6026 4 3 2 5994 5991 
2 6027 1 6026  
2 6028 1 6026  
2 6029 1 6026  
0 6030 4 1 2 5961 5997 
0 6031 4 1 2 5998 5958 
0 6032 4 2 2 6000 6001 
2 6033 1 6032  
2 6034 1 6032  
0 6035 4 1 2 5974 6006 
0 6036 4 1 2 6007 5932 
0 6037 4 2 2 6009 6010 
2 6038 1 6037  
2 6039 1 6037  
0 6040 4 3 2 6012 685 
2 6041 1 6040  
2 6042 1 6040  
2 6043 1 6040  
0 6044 4 1 2 5983 6015 
0 6045 4 1 2 6016 734 
0 6046 4 2 2 5901 6017 
2 6047 1 6046  
2 6048 1 6046  
0 6049 4 2 2 6018 6019 
2 6050 1 6049  
2 6051 1 6049  
0 6052 4 3 2 6024 6021 
2 6053 1 6052  
2 6054 1 6052  
2 6055 1 6052  
0 6056 4 1 2 5995 6027 
0 6057 4 1 2 6028 5992 
0 6058 4 2 2 6030 6031 
2 6059 1 6058  
2 6060 1 6058  
0 6061 4 2 2 6035 6036 
2 6062 1 6061  
2 6063 1 6061  
0 6064 4 3 2 6038 637 
2 6065 1 6064  
2 6066 1 6064  
2 6067 1 6064  
0 6068 4 1 2 6013 6041 
0 6069 4 1 2 6042 686 
0 6070 4 2 2 5944 6043 
2 6071 1 6070  
2 6072 1 6070  
0 6073 4 2 2 6044 6045 
2 6074 1 6073  
2 6075 1 6073  
0 6076 4 3 2 6050 6047 
2 6077 1 6076  
2 6078 1 6076  
2 6079 1 6076  
0 6080 4 1 2 6025 6053 
0 6081 4 1 2 6054 6022 
0 6082 4 2 2 6056 6057 
2 6083 1 6082  
2 6084 1 6082  
0 6085 4 3 2 6062 589 
2 6086 1 6085  
2 6087 1 6085  
2 6088 1 6085  
0 6089 4 1 2 6039 6065 
0 6090 4 1 2 6066 638 
0 6091 4 2 2 5978 6067 
2 6092 1 6091  
2 6093 1 6091  
0 6094 4 2 2 6068 6069 
2 6095 1 6094  
2 6096 1 6094  
0 6097 4 3 2 6074 6071 
2 6098 1 6097  
2 6099 1 6097  
2 6100 1 6097  
0 6101 4 1 2 6051 6077 
0 6102 4 1 2 6078 6048 
0 6103 4 2 2 6080 6081 
2 6104 1 6103  
2 6105 1 6103  
0 6106 4 1 2 6063 6086 
0 6107 4 1 2 6087 590 
0 6108 4 2 2 6008 6088 
2 6109 1 6108  
2 6110 1 6108  
0 6111 4 2 2 6089 6090 
2 6112 1 6111  
2 6113 1 6111  
0 6114 4 3 2 6095 6092 
2 6115 1 6114  
2 6116 1 6114  
2 6117 1 6114  
0 6118 4 1 2 6075 6098 
0 6119 4 1 2 6099 6072 
0 6120 4 2 2 6101 6102 
2 6121 1 6120  
2 6122 1 6120  
3 6123 4 0 2 6106 6107 
0 6124 4 3 2 6112 6109 
2 6125 1 6124  
2 6126 1 6124  
2 6127 1 6124  
0 6128 4 1 2 6096 6115 
0 6129 4 1 2 6116 6093 
0 6130 4 2 2 6118 6119 
2 6131 1 6130  
2 6132 1 6130  
0 6133 4 1 2 6113 6125 
0 6134 4 1 2 6126 6110 
0 6135 4 2 2 6128 6129 
2 6136 1 6135  
2 6137 1 6135  
0 6138 4 2 2 6133 6134 
2 6139 1 6138  
2 6140 1 6138  
0 6141 5 3 1 6139 
2 6142 1 6141  
2 6143 1 6141  
2 6144 1 6141  
0 6145 4 1 2 6140 6142 
0 6146 5 1 1 6143 
0 6147 4 2 2 6127 6144 
2 6148 1 6147  
2 6149 1 6147  
3 6150 4 0 2 6145 6146 
0 6151 4 3 2 6136 6148 
2 6152 1 6151  
2 6153 1 6151  
2 6154 1 6151  
0 6155 4 1 2 6137 6152 
0 6156 4 1 2 6153 6149 
0 6157 4 2 2 6117 6154 
2 6158 1 6157  
2 6159 1 6157  
3 6160 4 0 2 6155 6156 
0 6161 4 3 2 6131 6158 
2 6162 1 6161  
2 6163 1 6161  
2 6164 1 6161  
0 6165 4 1 2 6132 6162 
0 6166 4 1 2 6163 6159 
0 6167 4 2 2 6100 6164 
2 6168 1 6167  
2 6169 1 6167  
3 6170 4 0 2 6165 6166 
0 6171 4 3 2 6121 6168 
2 6172 1 6171  
2 6173 1 6171  
2 6174 1 6171  
0 6175 4 1 2 6122 6172 
0 6176 4 1 2 6173 6169 
0 6177 4 2 2 6079 6174 
2 6178 1 6177  
2 6179 1 6177  
3 6180 4 0 2 6175 6176 
0 6181 4 3 2 6104 6178 
2 6182 1 6181  
2 6183 1 6181  
2 6184 1 6181  
0 6185 4 1 2 6105 6182 
0 6186 4 1 2 6183 6179 
0 6187 4 2 2 6055 6184 
2 6188 1 6187  
2 6189 1 6187  
3 6190 4 0 2 6185 6186 
0 6191 4 3 2 6083 6188 
2 6192 1 6191  
2 6193 1 6191  
2 6194 1 6191  
0 6195 4 1 2 6084 6192 
0 6196 4 1 2 6193 6189 
0 6197 4 2 2 6029 6194 
2 6198 1 6197  
2 6199 1 6197  
3 6200 4 0 2 6195 6196 
0 6201 4 3 2 6059 6198 
2 6202 1 6201  
2 6203 1 6201  
2 6204 1 6201  
0 6205 4 1 2 6060 6202 
0 6206 4 1 2 6203 6199 
0 6207 4 2 2 5999 6204 
2 6208 1 6207  
2 6209 1 6207  
3 6210 4 0 2 6205 6206 
0 6211 4 3 2 6033 6208 
2 6212 1 6211  
2 6213 1 6211  
2 6214 1 6211  
0 6215 4 1 2 6034 6212 
0 6216 4 1 2 6213 6209 
0 6217 4 2 2 5965 6214 
2 6218 1 6217  
2 6219 1 6217  
3 6220 4 0 2 6215 6216 
0 6221 4 3 2 6003 6218 
2 6222 1 6221  
2 6223 1 6221  
2 6224 1 6221  
0 6225 4 1 2 6004 6222 
0 6226 4 1 2 6223 6219 
0 6227 4 2 2 5922 6224 
2 6228 1 6227  
2 6229 1 6227  
3 6230 4 0 2 6225 6226 
0 6231 4 3 2 5969 6228 
2 6232 1 6231  
2 6233 1 6231  
2 6234 1 6231  
0 6235 4 1 2 5970 6232 
0 6236 4 1 2 6233 6229 
0 6237 4 2 2 5876 6234 
2 6238 1 6237  
2 6239 1 6237  
3 6240 4 0 2 6235 6236 
0 6241 4 3 2 5926 6238 
2 6242 1 6241  
2 6243 1 6241  
2 6244 1 6241  
0 6245 4 1 2 5927 6242 
0 6246 4 1 2 6243 6239 
0 6247 4 2 2 5828 6244 
2 6248 1 6247  
2 6249 1 6247  
3 6250 4 0 2 6245 6246 
0 6251 4 3 2 5880 6248 
2 6252 1 6251  
2 6253 1 6251  
2 6254 1 6251  
0 6255 4 1 2 5881 6252 
0 6256 4 1 2 6253 6249 
0 6257 4 2 2 5779 6254 
2 6258 1 6257  
2 6259 1 6257  
3 6260 4 0 2 6255 6256 
0 6261 4 3 2 5832 6258 
2 6262 1 6261  
2 6263 1 6261  
2 6264 1 6261  
0 6265 4 1 2 5833 6262 
0 6266 4 1 2 6263 6259 
0 6267 4 2 2 5724 6264 
2 6268 1 6267  
2 6269 1 6267  
3 6270 4 0 2 6265 6266 
0 6271 4 3 2 5783 6268 
2 6272 1 6271  
2 6273 1 6271  
2 6274 1 6271  
0 6275 4 1 2 5784 6272 
0 6276 4 1 2 6273 6269 
0 6277 4 2 2 5669 6274 
2 6278 1 6277  
2 6279 1 6277  
3 6280 4 0 2 6275 6276 
0 6281 4 3 2 5728 6278 
2 6282 1 6281  
2 6283 1 6281  
2 6284 1 6281  
0 6285 4 1 2 5729 6282 
0 6286 4 1 2 6283 6279 
3 6287 4 0 2 5605 6284 
3 6288 4 0 2 6285 6286 
