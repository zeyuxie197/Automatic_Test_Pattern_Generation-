1 1 0 3 0 
2 2 1 1  
2 3 1 1  
2 4 1 1  
1 5 0 3 0 
2 6 1 5  
2 7 1 5  
2 8 1 5  
1 9 0 3 0 
2 10 1 9  
2 11 1 9  
2 12 1 9  
1 13 0 3 0 
2 14 1 13  
2 15 1 13  
2 16 1 13  
1 17 0 3 0 
2 18 1 17  
2 19 1 17  
2 20 1 17  
1 21 0 3 0 
2 22 1 21  
2 23 1 21  
2 24 1 21  
1 25 0 3 0 
2 26 1 25  
2 27 1 25  
2 28 1 25  
1 29 0 3 0 
2 30 1 29  
2 31 1 29  
2 32 1 29  
1 33 0 3 0 
2 34 1 33  
2 35 1 33  
2 36 1 33  
1 37 0 3 0 
2 38 1 37  
2 39 1 37  
2 40 1 37  
1 41 0 3 0 
2 42 1 41  
2 43 1 41  
2 44 1 41  
0 554 5 1 1 355 
0 555 5 1 1 368 
0 556 5 1 1 381 
1 45 0 3 0 
2 46 1 45  
2 47 1 45  
2 48 1 45  
0 557 5 1 1 356 
0 558 5 1 1 369 
0 559 5 1 1 394 
1 49 0 3 0 
2 50 1 49  
2 51 1 49  
2 52 1 49  
0 560 5 1 1 357 
0 561 5 1 1 382 
0 562 5 1 1 395 
1 53 0 3 0 
2 54 1 53  
2 55 1 53  
2 56 1 53  
0 563 5 1 1 370 
0 564 5 1 1 383 
0 565 5 1 1 396 
1 57 0 3 0 
2 58 1 57  
2 59 1 57  
2 60 1 57  
0 566 5 1 1 420 
0 567 5 1 1 446 
0 568 5 1 1 421 
1 61 0 3 0 
2 62 1 61  
2 63 1 61  
2 64 1 61  
0 569 5 1 1 433 
0 570 5 1 1 407 
0 571 5 1 1 447 
1 65 0 3 0 
2 66 1 65  
2 67 1 65  
2 68 1 65  
0 572 5 1 1 408 
0 573 5 1 1 434 
0 574 5 1 1 409 
1 69 0 3 0 
2 70 1 69  
2 71 1 69  
2 72 1 69  
0 575 5 1 1 422 
0 576 5 1 1 435 
0 577 5 1 1 410 
1 73 0 3 0 
2 74 1 73  
2 75 1 73  
2 76 1 73  
0 578 5 1 1 423 
0 579 5 1 1 448 
0 580 5 1 1 411 
1 77 0 3 0 
2 78 1 77  
2 79 1 77  
2 80 1 77  
0 581 5 1 1 436 
0 582 5 1 1 449 
0 583 5 1 1 424 
1 81 0 3 0 
2 82 1 81  
2 83 1 81  
2 84 1 81  
0 585 5 1 1 450 
0 586 5 1 1 371 
0 587 5 1 1 397 
1 85 0 3 0 
2 86 1 85  
2 87 1 85  
2 88 1 85  
0 589 5 1 1 384 
0 590 5 1 1 358 
0 591 5 1 1 398 
1 89 0 3 0 
2 90 1 89  
2 91 1 89  
2 92 1 89  
0 593 5 1 1 385 
0 594 7 1 4 554 555 556 399 
0 595 7 1 4 557 558 386 559 
1 93 0 3 0 
2 94 1 93  
2 95 1 93  
2 96 1 93  
0 597 7 1 4 360 563 564 565 
0 598 7 1 4 574 575 576 451 
0 599 7 1 4 577 578 438 579 
1 97 0 3 0 
2 98 1 97  
2 99 1 97  
2 100 1 97  
0 601 7 1 4 412 583 584 585 
0 602 3 4 4 594 595 596 597 
2 603 1 602  
2 604 1 602  
2 605 1 602  
2 606 1 602  
0 607 3 4 4 598 599 600 601 
2 608 1 607  
2 609 1 607  
2 610 1 607  
2 611 1 607  
1 101 0 3 0 
2 102 1 101  
2 103 1 101  
2 104 1 101  
1 105 0 3 0 
2 106 1 105  
2 107 1 105  
2 108 1 105  
0 620 7 4 5 413 566 439 567 603 
2 621 1 620  
2 622 1 620  
2 623 1 620  
2 624 1 620  
1 109 0 3 0 
2 110 1 109  
2 111 1 109  
2 112 1 109  
1 113 0 3 0 
2 114 1 113  
2 115 1 113  
2 116 1 113  
0 625 7 4 5 414 568 569 452 604 
2 626 1 625  
2 627 1 625  
2 628 1 625  
2 629 1 625  
1 117 0 3 0 
2 118 1 117  
2 119 1 117  
2 120 1 117  
0 630 7 4 5 570 426 440 571 605 
2 631 1 630  
2 632 1 630  
2 633 1 630  
2 634 1 630  
1 121 0 3 0 
2 122 1 121  
2 123 1 121  
2 124 1 121  
0 635 7 4 5 572 427 573 453 606 
2 636 1 635  
2 637 1 635  
2 638 1 635  
2 639 1 635  
1 125 0 3 0 
2 126 1 125  
2 127 1 125  
2 128 1 125  
0 640 7 4 5 361 586 387 587 608 
2 641 1 640  
2 642 1 640  
2 643 1 640  
2 644 1 640  
1 129 0 1 0 
1 130 0 1 0 
1 131 0 1 0 
1 132 0 1 0 
1 133 0 1 0 
1 134 0 1 0 
1 135 0 1 0 
1 136 0 1 0 
1 137 0 8 0 
2 138 1 137  
2 139 1 137  
2 140 1 137  
2 141 1 137  
2 142 1 137  
2 143 1 137  
2 144 1 137  
2 145 1 137  
0 645 7 4 5 362 588 589 400 609 
2 646 1 645  
2 647 1 645  
2 648 1 645  
2 649 1 645  
0 650 7 4 5 590 374 388 591 610 
2 651 1 650  
2 652 1 650  
2 653 1 650  
2 654 1 650  
0 655 7 4 5 592 375 593 401 611 
2 656 1 655  
2 657 1 655  
2 658 1 655  
2 659 1 655  
0 692 7 1 2 363 621 
0 693 7 1 2 376 622 
0 694 7 1 2 389 623 
0 695 7 1 2 402 624 
0 696 7 1 2 364 626 
0 697 7 1 2 377 627 
0 698 7 1 2 390 628 
0 699 7 1 2 403 629 
0 700 7 1 2 365 631 
0 701 7 1 2 378 632 
0 702 7 1 2 391 633 
0 703 7 1 2 404 634 
0 704 7 1 2 366 636 
0 705 7 1 2 379 637 
0 706 7 1 2 392 638 
0 707 7 1 2 405 639 
0 708 7 1 2 415 641 
0 709 7 1 2 428 642 
0 710 7 1 2 441 643 
0 711 7 1 2 454 644 
0 712 7 1 2 416 646 
0 713 7 1 2 429 647 
0 714 7 1 2 442 648 
0 715 7 1 2 455 649 
0 716 7 1 2 417 651 
0 717 7 1 2 430 652 
0 718 7 1 2 443 653 
0 719 7 1 2 456 654 
0 720 7 1 2 418 656 
0 721 7 1 2 431 657 
0 722 7 1 2 444 658 
0 723 7 1 2 457 659 
3 724 2 0 2 4 692 
3 725 2 0 2 8 693 
3 726 2 0 2 12 694 
3 727 2 0 2 16 695 
3 728 2 0 2 20 696 
3 729 2 0 2 24 697 
3 730 2 0 2 28 698 
3 731 2 0 2 32 699 
3 732 2 0 2 36 700 
3 733 2 0 2 40 701 
3 734 2 0 2 44 702 
3 735 2 0 2 48 703 
3 736 2 0 2 52 704 
3 737 2 0 2 56 705 
3 738 2 0 2 60 706 
3 739 2 0 2 64 707 
3 740 2 0 2 68 708 
3 741 2 0 2 72 709 
3 742 2 0 2 76 710 
3 743 2 0 2 80 711 
3 744 2 0 2 84 712 
3 745 2 0 2 88 713 
3 746 2 0 2 92 714 
3 747 2 0 2 96 715 
3 748 2 0 2 100 716 
3 749 2 0 2 104 717 
3 750 2 0 2 108 718 
3 751 2 0 2 112 719 
3 752 2 0 2 116 720 
3 753 2 0 2 120 721 
3 754 2 0 2 124 722 
3 755 2 0 2 128 723 
0 250 2 1 2 2 6 
0 251 2 1 2 10 14 
0 252 2 1 2 18 22 
0 253 2 1 2 26 30 
0 254 2 1 2 34 38 
0 255 2 1 2 42 46 
0 256 2 1 2 50 54 
0 257 2 1 2 58 62 
0 258 2 1 2 66 70 
0 259 2 1 2 74 78 
0 260 2 1 2 82 86 
0 261 2 1 2 90 94 
0 262 2 1 2 98 102 
0 263 2 1 2 106 110 
0 264 2 1 2 114 118 
0 265 2 1 2 122 126 
0 266 7 1 2 129 138 
0 267 7 1 2 130 139 
0 268 7 1 2 131 140 
0 269 7 1 2 132 141 
0 270 7 1 2 133 142 
0 271 7 1 2 134 143 
0 272 7 1 2 135 144 
0 273 7 1 2 136 145 
0 274 2 1 2 3 19 
0 275 2 1 2 35 51 
0 276 2 1 2 7 23 
0 277 2 1 2 39 55 
0 278 2 1 2 11 27 
0 279 2 1 2 43 59 
0 280 2 1 2 15 31 
0 281 2 1 2 47 63 
0 282 2 1 2 67 83 
0 283 2 1 2 99 115 
0 284 2 1 2 71 87 
0 285 2 1 2 103 119 
0 286 2 1 2 75 91 
0 287 2 1 2 107 123 
0 288 2 1 2 79 95 
0 289 2 1 2 111 127 
0 290 2 2 2 250 251 
2 291 1 290  
2 292 1 290  
0 293 2 2 2 252 253 
2 294 1 293  
2 295 1 293  
0 296 2 2 2 254 255 
2 297 1 296  
2 298 1 296  
0 299 2 2 2 256 257 
2 300 1 299  
2 301 1 299  
0 302 2 2 2 258 259 
2 303 1 302  
2 304 1 302  
0 305 2 2 2 260 261 
2 306 1 305  
2 307 1 305  
0 308 2 2 2 262 263 
2 309 1 308  
2 310 1 308  
0 311 2 2 2 264 265 
2 312 1 311  
2 313 1 311  
0 314 2 1 2 274 275 
0 315 2 1 2 276 277 
0 316 2 1 2 278 279 
0 317 2 1 2 280 281 
0 318 2 1 2 282 283 
0 319 2 1 2 284 285 
0 320 2 1 2 286 287 
0 321 2 1 2 288 289 
0 338 2 1 2 291 294 
0 339 2 1 2 297 300 
0 340 2 1 2 292 298 
0 341 2 1 2 295 301 
0 342 2 1 2 303 306 
0 343 2 1 2 309 312 
0 344 2 1 2 304 310 
0 345 2 1 2 307 313 
0 346 2 1 2 266 342 
0 347 2 1 2 267 343 
0 348 2 1 2 268 344 
0 349 2 1 2 269 345 
0 350 2 1 2 270 338 
0 351 2 1 2 271 339 
0 352 2 1 2 272 340 
0 353 2 1 2 273 341 
0 354 2 12 2 314 346 
2 355 1 354  
2 356 1 354  
2 357 1 354  
2 358 1 354  
2 359 1 354  
2 360 1 354  
2 361 1 354  
2 362 1 354  
2 363 1 354  
2 364 1 354  
2 365 1 354  
2 366 1 354  
0 367 2 12 2 315 347 
2 368 1 367  
2 369 1 367  
2 370 1 367  
2 371 1 367  
2 372 1 367  
2 373 1 367  
2 374 1 367  
2 375 1 367  
2 376 1 367  
2 377 1 367  
2 378 1 367  
2 379 1 367  
0 584 5 1 1 437 
0 380 2 12 2 316 348 
2 381 1 380  
2 382 1 380  
2 383 1 380  
2 384 1 380  
2 385 1 380  
2 386 1 380  
2 387 1 380  
2 388 1 380  
2 389 1 380  
2 390 1 380  
2 391 1 380  
2 392 1 380  
0 393 2 12 2 317 349 
2 394 1 393  
2 395 1 393  
2 396 1 393  
2 397 1 393  
2 398 1 393  
2 399 1 393  
2 400 1 393  
2 401 1 393  
2 402 1 393  
2 403 1 393  
2 404 1 393  
2 405 1 393  
0 588 5 1 1 372 
0 406 2 12 2 318 350 
2 407 1 406  
2 408 1 406  
2 409 1 406  
2 410 1 406  
2 411 1 406  
2 412 1 406  
2 413 1 406  
2 414 1 406  
2 415 1 406  
2 416 1 406  
2 417 1 406  
2 418 1 406  
0 419 2 12 2 319 351 
2 420 1 419  
2 421 1 419  
2 422 1 419  
2 423 1 419  
2 424 1 419  
2 425 1 419  
2 426 1 419  
2 427 1 419  
2 428 1 419  
2 429 1 419  
2 430 1 419  
2 431 1 419  
0 592 5 1 1 359 
0 432 2 12 2 320 352 
2 433 1 432  
2 434 1 432  
2 435 1 432  
2 436 1 432  
2 437 1 432  
2 438 1 432  
2 439 1 432  
2 440 1 432  
2 441 1 432  
2 442 1 432  
2 443 1 432  
2 444 1 432  
0 596 7 1 4 560 373 561 562 
0 445 2 12 2 321 353 
2 446 1 445  
2 447 1 445  
2 448 1 445  
2 449 1 445  
2 450 1 445  
2 451 1 445  
2 452 1 445  
2 453 1 445  
2 454 1 445  
2 455 1 445  
2 456 1 445  
2 457 1 445  
0 600 7 1 4 580 425 581 582 
