1 0 0 6 0
1 1 0 6 0
1 2 0 6 0
1 3 0 6 0
1 4 0 6 0
1 5 0 6 0
1 6 0 6 0
1 7 0 6 0
1 8 0 6 0
1 9 0 6 0
1 10 0 6 0
1 11 0 6 0
1 12 0 6 0
1 13 0 6 0
1 14 0 6 0
1 15 0 6 0
1 16 0 6 0
1 17 0 6 0
1 18 0 6 0
1 19 0 6 0
1 20 0 6 0
1 21 0 6 0
1 22 0 6 0
1 23 0 6 0
1 24 0 6 0
1 25 0 6 0
1 26 0 6 0
1 27 0 6 0
1 28 0 6 0
1 29 0 6 0
1 30 0 6 0
1 31 0 6 0
1 32 0 1 0
1 33 0 1 0
1 34 0 1 0
1 35 0 1 0
1 36 0 1 0
1 37 0 1 0
1 38 0 1 0
1 39 0 1 0
1 40 0 8 0
3 41 5 0 1 555 
3 42 5 0 1 556 
3 43 5 0 1 557 
3 44 5 0 1 558 
3 45 5 0 1 559 
3 46 5 0 1 560 
3 47 5 0 1 561 
3 48 5 0 1 562 
3 49 5 0 1 563 
3 50 5 0 1 564 
3 51 5 0 1 565 
3 52 5 0 1 566 
3 53 5 0 1 567 
3 54 5 0 1 568 
3 55 5 0 1 569 
3 56 5 0 1 570 
3 57 5 0 1 571 
3 58 5 0 1 572 
3 59 5 0 1 573 
3 60 5 0 1 574 
3 61 5 0 1 575 
3 62 5 0 1 576 
3 63 5 0 1 577 
3 64 5 0 1 578 
3 65 5 0 1 579 
3 66 5 0 1 580 
3 67 5 0 1 581 
3 68 5 0 1 582 
3 69 5 0 1 583 
3 70 5 0 1 584 
3 71 5 0 1 585 
3 72 5 0 1 586 
0 73 7 2 2 32 779 
0 74 7 2 2 33 780 
0 75 7 2 2 34 781 
0 76 7 2 2 35 782 
0 77 7 2 2 36 783 
0 78 7 2 2 37 784 
0 79 7 2 2 38 785 
0 80 7 2 2 39 786 
0 81 6 2 2 587 593 
0 82 6 2 2 599 605 
0 83 6 2 2 611 617 
0 84 6 2 2 623 629 
0 85 6 2 2 635 641 
0 86 6 2 2 647 653 
0 87 6 2 2 659 665 
0 88 6 2 2 671 677 
0 89 6 2 2 683 689 
0 90 6 2 2 695 701 
0 91 6 2 2 707 713 
0 92 6 2 2 719 725 
0 93 6 2 2 731 737 
0 94 6 2 2 743 749 
0 95 6 2 2 755 761 
0 96 6 2 2 767 773 
0 97 6 2 2 588 612 
0 98 6 2 2 636 660 
0 99 6 2 2 594 618 
0 100 6 2 2 642 666 
0 101 6 2 2 600 624 
0 102 6 2 2 648 672 
0 103 6 2 2 606 630 
0 104 6 2 2 654 678 
0 105 6 2 2 684 708 
0 106 6 2 2 732 756 
0 107 6 2 2 690 714 
0 108 6 2 2 738 762 
0 109 6 2 2 696 720 
0 110 6 2 2 744 768 
0 111 6 2 2 702 726 
0 112 6 2 2 750 774 
0 113 6 1 2 589 803 
0 114 6 1 2 595 804 
0 115 6 1 2 601 805 
0 116 6 1 2 607 806 
0 117 6 1 2 613 807 
0 118 6 1 2 619 808 
0 119 6 1 2 625 809 
0 120 6 1 2 631 810 
0 121 6 1 2 637 811 
0 122 6 1 2 643 812 
0 123 6 1 2 649 813 
0 124 6 1 2 655 814 
0 125 6 1 2 661 815 
0 126 6 1 2 667 816 
0 127 6 1 2 673 817 
0 128 6 1 2 679 818 
0 129 6 1 2 685 819 
0 130 6 1 2 691 820 
0 131 6 1 2 697 821 
0 132 6 1 2 703 822 
0 133 6 1 2 709 823 
0 134 6 1 2 715 824 
0 135 6 1 2 721 825 
0 136 6 1 2 727 826 
0 137 6 1 2 733 827 
0 138 6 1 2 739 828 
0 139 6 1 2 745 829 
0 140 6 1 2 751 830 
0 141 6 1 2 757 831 
0 142 6 1 2 763 832 
0 143 6 1 2 769 833 
0 144 6 1 2 775 834 
0 145 6 1 2 590 835 
0 146 6 1 2 614 836 
0 147 6 1 2 638 837 
0 148 6 1 2 662 838 
0 149 6 1 2 596 839 
0 150 6 1 2 620 840 
0 151 6 1 2 644 841 
0 152 6 1 2 668 842 
0 153 6 1 2 602 843 
0 154 6 1 2 626 844 
0 155 6 1 2 650 845 
0 156 6 1 2 674 846 
0 157 6 1 2 608 847 
0 158 6 1 2 632 848 
0 159 6 1 2 656 849 
0 160 6 1 2 680 850 
0 161 6 1 2 686 851 
0 162 6 1 2 710 852 
0 163 6 1 2 734 853 
0 164 6 1 2 758 854 
0 165 6 1 2 692 855 
0 166 6 1 2 716 856 
0 167 6 1 2 740 857 
0 168 6 1 2 764 858 
0 169 6 1 2 698 859 
0 170 6 1 2 722 860 
0 171 6 1 2 746 861 
0 172 6 1 2 770 862 
0 173 6 1 2 704 863 
0 174 6 1 2 728 864 
0 175 6 1 2 752 865 
0 176 6 1 2 776 866 
0 177 6 2 2 113 114 
0 178 6 2 2 115 116 
0 179 6 2 2 117 118 
0 180 6 2 2 119 120 
0 181 6 2 2 121 122 
0 182 6 2 2 123 124 
0 183 6 2 2 125 126 
0 184 6 2 2 127 128 
0 185 6 2 2 129 130 
0 186 6 2 2 131 132 
0 187 6 2 2 133 134 
0 188 6 2 2 135 136 
0 189 6 2 2 137 138 
0 190 6 2 2 139 140 
0 191 6 2 2 141 142 
0 192 6 2 2 143 144 
0 193 6 2 2 145 146 
0 194 6 2 2 147 148 
0 195 6 2 2 149 150 
0 196 6 2 2 151 152 
0 197 6 2 2 153 154 
0 198 6 2 2 155 156 
0 199 6 2 2 157 158 
0 200 6 2 2 159 160 
0 201 6 2 2 161 162 
0 202 6 2 2 163 164 
0 203 6 2 2 165 166 
0 204 6 2 2 167 168 
0 205 6 2 2 169 170 
0 206 6 2 2 171 172 
0 207 6 2 2 173 174 
0 208 6 2 2 175 176 
0 209 6 2 2 867 869 
0 210 6 2 2 871 873 
0 211 6 2 2 875 877 
0 212 6 2 2 879 881 
0 213 6 2 2 883 885 
0 214 6 2 2 887 889 
0 215 6 2 2 891 893 
0 216 6 2 2 895 897 
0 217 6 2 2 899 901 
0 218 6 2 2 903 905 
0 219 6 2 2 907 909 
0 220 6 2 2 911 913 
0 221 6 2 2 915 917 
0 222 6 2 2 919 921 
0 223 6 2 2 923 925 
0 224 6 2 2 927 929 
0 225 6 1 2 868 931 
0 226 6 1 2 870 932 
0 227 6 1 2 872 933 
0 228 6 1 2 874 934 
0 229 6 1 2 876 935 
0 230 6 1 2 878 936 
0 231 6 1 2 880 937 
0 232 6 1 2 882 938 
0 233 6 1 2 884 939 
0 234 6 1 2 886 940 
0 235 6 1 2 888 941 
0 236 6 1 2 890 942 
0 237 6 1 2 892 943 
0 238 6 1 2 894 944 
0 239 6 1 2 896 945 
0 240 6 1 2 898 946 
0 241 6 1 2 900 947 
0 242 6 1 2 902 948 
0 243 6 1 2 904 949 
0 244 6 1 2 906 950 
0 245 6 1 2 908 951 
0 246 6 1 2 910 952 
0 247 6 1 2 912 953 
0 248 6 1 2 914 954 
0 249 6 1 2 916 955 
0 250 6 1 2 918 956 
0 251 6 1 2 920 957 
0 252 6 1 2 922 958 
0 253 6 1 2 924 959 
0 254 6 1 2 926 960 
0 255 6 1 2 928 961 
0 256 6 1 2 930 962 
0 257 6 4 2 225 226 
0 258 6 4 2 227 228 
0 259 6 4 2 229 230 
0 260 6 4 2 231 232 
0 261 6 4 2 233 234 
0 262 6 4 2 235 236 
0 263 6 4 2 237 238 
0 264 6 4 2 239 240 
0 265 6 2 2 241 242 
0 266 6 2 2 243 244 
0 267 6 2 2 245 246 
0 268 6 2 2 247 248 
0 269 6 2 2 249 250 
0 270 6 2 2 251 252 
0 271 6 2 2 253 254 
0 272 6 2 2 255 256 
0 273 6 2 2 963 967 
0 274 6 2 2 971 975 
0 275 6 2 2 964 972 
0 276 6 2 2 968 976 
0 277 6 2 2 979 983 
0 278 6 2 2 987 991 
0 279 6 2 2 980 988 
0 280 6 2 2 984 992 
0 281 6 1 2 965 1011 
0 282 6 1 2 969 1012 
0 283 6 1 2 973 1013 
0 284 6 1 2 977 1014 
0 285 6 1 2 966 1015 
0 286 6 1 2 974 1016 
0 287 6 1 2 970 1017 
0 288 6 1 2 978 1018 
0 289 6 1 2 981 1019 
0 290 6 1 2 985 1020 
0 291 6 1 2 989 1021 
0 292 6 1 2 993 1022 
0 293 6 1 2 982 1023 
0 294 6 1 2 990 1024 
0 295 6 1 2 986 1025 
0 296 6 1 2 994 1026 
0 297 6 2 2 281 282 
0 298 6 2 2 283 284 
0 299 6 2 2 285 286 
0 300 6 2 2 287 288 
0 301 6 2 2 289 290 
0 302 6 2 2 291 292 
0 303 6 2 2 293 294 
0 304 6 2 2 295 296 
0 305 6 2 2 787 1035 
0 306 6 2 2 789 1037 
0 307 6 2 2 791 1039 
0 308 6 2 2 793 1041 
0 309 6 2 2 795 1027 
0 310 6 2 2 797 1029 
0 311 6 2 2 799 1031 
0 312 6 2 2 801 1033 
0 313 6 1 2 788 1043 
0 314 6 1 2 1036 1044 
0 315 6 1 2 790 1045 
0 316 6 1 2 1038 1046 
0 317 6 1 2 792 1047 
0 318 6 1 2 1040 1048 
0 319 6 1 2 794 1049 
0 320 6 1 2 1042 1050 
0 321 6 1 2 796 1051 
0 322 6 1 2 1028 1052 
0 323 6 1 2 798 1053 
0 324 6 1 2 1030 1054 
0 325 6 1 2 800 1055 
0 326 6 1 2 1032 1056 
0 327 6 1 2 802 1057 
0 328 6 1 2 1034 1058 
0 329 6 2 2 313 314 
0 330 6 2 2 315 316 
0 331 6 2 2 317 318 
0 332 6 2 2 319 320 
0 333 6 2 2 321 322 
0 334 6 2 2 323 324 
0 335 6 2 2 325 326 
0 336 6 2 2 327 328 
0 337 6 2 2 995 1059 
0 338 6 2 2 997 1061 
0 339 6 2 2 999 1063 
0 340 6 2 2 1001 1065 
0 341 6 2 2 1003 1067 
0 342 6 2 2 1005 1069 
0 343 6 2 2 1007 1071 
0 344 6 2 2 1009 1073 
0 345 6 1 2 996 1075 
0 346 6 1 2 1060 1076 
0 347 6 1 2 998 1077 
0 348 6 1 2 1062 1078 
0 349 6 1 2 1000 1079 
0 350 6 1 2 1064 1080 
0 351 6 1 2 1002 1081 
0 352 6 1 2 1066 1082 
0 353 6 1 2 1004 1083 
0 354 6 1 2 1068 1084 
0 355 6 1 2 1006 1085 
0 356 6 1 2 1070 1086 
0 357 6 1 2 1008 1087 
0 358 6 1 2 1072 1088 
0 359 6 1 2 1010 1089 
0 360 6 1 2 1074 1090 
0 361 6 12 2 345 346 
0 362 6 12 2 347 348 
0 363 6 12 2 349 350 
0 364 6 12 2 351 352 
0 365 6 12 2 355 356 
0 366 6 12 2 359 360 
0 367 6 12 2 357 358 
0 368 6 12 2 353 354 
0 369 5 1 1 1091 
0 370 5 1 1 1103 
0 371 5 1 1 1115 
0 372 5 1 1 1092 
0 373 5 1 1 1104 
0 374 5 1 1 1127 
0 375 5 1 1 1093 
0 376 5 1 1 1116 
0 377 5 1 1 1128 
0 378 5 1 1 1105 
0 379 5 1 1 1117 
0 380 5 1 1 1129 
0 381 5 1 1 1139 
0 382 5 1 1 1151 
0 383 5 1 1 1140 
0 384 5 1 1 1163 
0 385 5 1 1 1175 
0 386 5 1 1 1152 
0 387 5 1 1 1176 
0 388 5 1 1 1164 
0 389 5 1 1 1177 
0 390 5 1 1 1141 
0 391 5 1 1 1165 
0 392 5 1 1 1178 
0 393 5 1 1 1142 
0 394 5 1 1 1153 
0 395 5 1 1 1179 
0 396 5 1 1 1166 
0 397 5 1 1 1154 
0 398 5 1 1 1143 
0 399 5 1 1 1167 
0 400 5 1 1 1155 
0 401 5 1 1 1106 
0 402 5 1 1 1130 
0 403 5 1 1 1107 
0 404 5 1 1 1118 
0 405 5 1 1 1094 
0 406 5 1 1 1131 
0 407 5 1 1 1095 
0 408 5 1 1 1119 
0 409 7 1 4 369 370 371 1132 
0 410 7 1 4 372 373 1120 374 
0 411 7 1 4 375 1108 376 377 
0 412 7 1 4 1096 378 379 380 
0 413 7 1 4 389 390 391 1156 
0 414 7 1 4 392 393 1168 394 
0 415 7 1 4 395 1144 396 397 
0 416 7 1 4 1180 398 399 400 
0 417 3 4 4 409 410 411 412 
0 418 3 4 4 413 414 415 416 
0 419 7 4 5 1181 381 1169 382 1187 
0 420 7 4 5 1182 383 384 1157 1188 
0 421 7 4 5 385 1145 1170 386 1189 
0 422 7 4 5 387 1146 388 1158 1190 
0 423 7 4 5 1097 401 1121 402 1191 
0 424 7 4 5 1098 403 404 1133 1192 
0 425 7 4 5 405 1109 1122 406 1193 
0 426 7 4 5 407 1110 408 1134 1194 
0 427 7 2 2 1099 1195 
0 428 7 2 2 1111 1196 
0 429 7 2 2 1123 1197 
0 430 7 2 2 1135 1198 
0 431 7 2 2 1100 1199 
0 432 7 2 2 1112 1200 
0 433 7 2 2 1124 1201 
0 434 7 2 2 1136 1202 
0 435 7 2 2 1101 1203 
0 436 7 2 2 1113 1204 
0 437 7 2 2 1125 1205 
0 438 7 2 2 1137 1206 
0 439 7 2 2 1102 1207 
0 440 7 2 2 1114 1208 
0 441 7 2 2 1126 1209 
0 442 7 2 2 1138 1210 
0 443 7 2 2 1183 1211 
0 444 7 2 2 1147 1212 
0 445 7 2 2 1171 1213 
0 446 7 2 2 1159 1214 
0 447 7 2 2 1184 1215 
0 448 7 2 2 1148 1216 
0 449 7 2 2 1172 1217 
0 450 7 2 2 1160 1218 
0 451 7 2 2 1185 1219 
0 452 7 2 2 1149 1220 
0 453 7 2 2 1173 1221 
0 454 7 2 2 1161 1222 
0 455 7 2 2 1186 1223 
0 456 7 2 2 1150 1224 
0 457 7 2 2 1174 1225 
0 458 7 2 2 1162 1226 
0 459 6 2 2 591 1227 
0 460 6 2 2 597 1229 
0 461 6 2 2 603 1231 
0 462 6 2 2 609 1233 
0 463 6 2 2 615 1235 
0 464 6 2 2 621 1237 
0 465 6 2 2 627 1239 
0 466 6 2 2 633 1241 
0 467 6 2 2 639 1243 
0 468 6 2 2 645 1245 
0 469 6 2 2 651 1247 
0 470 6 2 2 657 1249 
0 471 6 2 2 663 1251 
0 472 6 2 2 669 1253 
0 473 6 2 2 675 1255 
0 474 6 2 2 681 1257 
0 475 6 2 2 687 1259 
0 476 6 2 2 693 1261 
0 477 6 2 2 699 1263 
0 478 6 2 2 705 1265 
0 479 6 2 2 711 1267 
0 480 6 2 2 717 1269 
0 481 6 2 2 723 1271 
0 482 6 2 2 729 1273 
0 483 6 2 2 735 1275 
0 484 6 2 2 741 1277 
0 485 6 2 2 747 1279 
0 486 6 2 2 753 1281 
0 487 6 2 2 759 1283 
0 488 6 2 2 765 1285 
0 489 6 2 2 771 1287 
0 490 6 2 2 777 1289 
0 491 6 1 2 592 1291 
0 492 6 1 2 1228 1292 
0 493 6 1 2 598 1293 
0 494 6 1 2 1230 1294 
0 495 6 1 2 604 1295 
0 496 6 1 2 1232 1296 
0 497 6 1 2 610 1297 
0 498 6 1 2 1234 1298 
0 499 6 1 2 616 1299 
0 500 6 1 2 1236 1300 
0 501 6 1 2 622 1301 
0 502 6 1 2 1238 1302 
0 503 6 1 2 628 1303 
0 504 6 1 2 1240 1304 
0 505 6 1 2 634 1305 
0 506 6 1 2 1242 1306 
0 507 6 1 2 640 1307 
0 508 6 1 2 1244 1308 
0 509 6 1 2 646 1309 
0 510 6 1 2 1246 1310 
0 511 6 1 2 652 1311 
0 512 6 1 2 1248 1312 
0 513 6 1 2 658 1313 
0 514 6 1 2 1250 1314 
0 515 6 1 2 664 1315 
0 516 6 1 2 1252 1316 
0 517 6 1 2 670 1317 
0 518 6 1 2 1254 1318 
0 519 6 1 2 676 1319 
0 520 6 1 2 1256 1320 
0 521 6 1 2 682 1321 
0 522 6 1 2 1258 1322 
0 523 6 1 2 688 1323 
0 524 6 1 2 1260 1324 
0 525 6 1 2 694 1325 
0 526 6 1 2 1262 1326 
0 527 6 1 2 700 1327 
0 528 6 1 2 1264 1328 
0 529 6 1 2 706 1329 
0 530 6 1 2 1266 1330 
0 531 6 1 2 712 1331 
0 532 6 1 2 1268 1332 
0 533 6 1 2 718 1333 
0 534 6 1 2 1270 1334 
0 535 6 1 2 724 1335 
0 536 6 1 2 1272 1336 
0 537 6 1 2 730 1337 
0 538 6 1 2 1274 1338 
0 539 6 1 2 736 1339 
0 540 6 1 2 1276 1340 
0 541 6 1 2 742 1341 
0 542 6 1 2 1278 1342 
0 543 6 1 2 748 1343 
0 544 6 1 2 1280 1344 
0 545 6 1 2 754 1345 
0 546 6 1 2 1282 1346 
0 547 6 1 2 760 1347 
0 548 6 1 2 1284 1348 
0 549 6 1 2 766 1349 
0 550 6 1 2 1286 1350 
0 551 6 1 2 772 1351 
0 552 6 1 2 1288 1352 
0 553 6 1 2 778 1353 
0 554 6 1 2 1290 1354 
0 555 6 1 2 491 492 
0 556 6 1 2 493 494 
0 557 6 1 2 495 496 
0 558 6 1 2 497 498 
0 559 6 1 2 499 500 
0 560 6 1 2 501 502 
0 561 6 1 2 503 504 
0 562 6 1 2 505 506 
0 563 6 1 2 507 508 
0 564 6 1 2 509 510 
0 565 6 1 2 511 512 
0 566 6 1 2 513 514 
0 567 6 1 2 515 516 
0 568 6 1 2 517 518 
0 569 6 1 2 519 520 
0 570 6 1 2 521 522 
0 571 6 1 2 523 524 
0 572 6 1 2 525 526 
0 573 6 1 2 527 528 
0 574 6 1 2 529 530 
0 575 6 1 2 531 532 
0 576 6 1 2 533 534 
0 577 6 1 2 535 536 
0 578 6 1 2 537 538 
0 579 6 1 2 539 540 
0 580 6 1 2 541 542 
0 581 6 1 2 543 544 
0 582 6 1 2 545 546 
0 583 6 1 2 547 548 
0 584 6 1 2 549 550 
0 585 6 1 2 551 552 
0 586 6 1 2 553 554 
2 587 1 0
2 588 1 0
2 589 1 0
2 590 1 0
2 591 1 0
2 592 1 0
2 593 1 1
2 594 1 1
2 595 1 1
2 596 1 1
2 597 1 1
2 598 1 1
2 599 1 2
2 600 1 2
2 601 1 2
2 602 1 2
2 603 1 2
2 604 1 2
2 605 1 3
2 606 1 3
2 607 1 3
2 608 1 3
2 609 1 3
2 610 1 3
2 611 1 4
2 612 1 4
2 613 1 4
2 614 1 4
2 615 1 4
2 616 1 4
2 617 1 5
2 618 1 5
2 619 1 5
2 620 1 5
2 621 1 5
2 622 1 5
2 623 1 6
2 624 1 6
2 625 1 6
2 626 1 6
2 627 1 6
2 628 1 6
2 629 1 7
2 630 1 7
2 631 1 7
2 632 1 7
2 633 1 7
2 634 1 7
2 635 1 8
2 636 1 8
2 637 1 8
2 638 1 8
2 639 1 8
2 640 1 8
2 641 1 9
2 642 1 9
2 643 1 9
2 644 1 9
2 645 1 9
2 646 1 9
2 647 1 10
2 648 1 10
2 649 1 10
2 650 1 10
2 651 1 10
2 652 1 10
2 653 1 11
2 654 1 11
2 655 1 11
2 656 1 11
2 657 1 11
2 658 1 11
2 659 1 12
2 660 1 12
2 661 1 12
2 662 1 12
2 663 1 12
2 664 1 12
2 665 1 13
2 666 1 13
2 667 1 13
2 668 1 13
2 669 1 13
2 670 1 13
2 671 1 14
2 672 1 14
2 673 1 14
2 674 1 14
2 675 1 14
2 676 1 14
2 677 1 15
2 678 1 15
2 679 1 15
2 680 1 15
2 681 1 15
2 682 1 15
2 683 1 16
2 684 1 16
2 685 1 16
2 686 1 16
2 687 1 16
2 688 1 16
2 689 1 17
2 690 1 17
2 691 1 17
2 692 1 17
2 693 1 17
2 694 1 17
2 695 1 18
2 696 1 18
2 697 1 18
2 698 1 18
2 699 1 18
2 700 1 18
2 701 1 19
2 702 1 19
2 703 1 19
2 704 1 19
2 705 1 19
2 706 1 19
2 707 1 20
2 708 1 20
2 709 1 20
2 710 1 20
2 711 1 20
2 712 1 20
2 713 1 21
2 714 1 21
2 715 1 21
2 716 1 21
2 717 1 21
2 718 1 21
2 719 1 22
2 720 1 22
2 721 1 22
2 722 1 22
2 723 1 22
2 724 1 22
2 725 1 23
2 726 1 23
2 727 1 23
2 728 1 23
2 729 1 23
2 730 1 23
2 731 1 24
2 732 1 24
2 733 1 24
2 734 1 24
2 735 1 24
2 736 1 24
2 737 1 25
2 738 1 25
2 739 1 25
2 740 1 25
2 741 1 25
2 742 1 25
2 743 1 26
2 744 1 26
2 745 1 26
2 746 1 26
2 747 1 26
2 748 1 26
2 749 1 27
2 750 1 27
2 751 1 27
2 752 1 27
2 753 1 27
2 754 1 27
2 755 1 28
2 756 1 28
2 757 1 28
2 758 1 28
2 759 1 28
2 760 1 28
2 761 1 29
2 762 1 29
2 763 1 29
2 764 1 29
2 765 1 29
2 766 1 29
2 767 1 30
2 768 1 30
2 769 1 30
2 770 1 30
2 771 1 30
2 772 1 30
2 773 1 31
2 774 1 31
2 775 1 31
2 776 1 31
2 777 1 31
2 778 1 31
2 779 1 40
2 780 1 40
2 781 1 40
2 782 1 40
2 783 1 40
2 784 1 40
2 785 1 40
2 786 1 40
2 787 1 73
2 788 1 73
2 789 1 74
2 790 1 74
2 791 1 75
2 792 1 75
2 793 1 76
2 794 1 76
2 795 1 77
2 796 1 77
2 797 1 78
2 798 1 78
2 799 1 79
2 800 1 79
2 801 1 80
2 802 1 80
2 803 1 81
2 804 1 81
2 805 1 82
2 806 1 82
2 807 1 83
2 808 1 83
2 809 1 84
2 810 1 84
2 811 1 85
2 812 1 85
2 813 1 86
2 814 1 86
2 815 1 87
2 816 1 87
2 817 1 88
2 818 1 88
2 819 1 89
2 820 1 89
2 821 1 90
2 822 1 90
2 823 1 91
2 824 1 91
2 825 1 92
2 826 1 92
2 827 1 93
2 828 1 93
2 829 1 94
2 830 1 94
2 831 1 95
2 832 1 95
2 833 1 96
2 834 1 96
2 835 1 97
2 836 1 97
2 837 1 98
2 838 1 98
2 839 1 99
2 840 1 99
2 841 1 100
2 842 1 100
2 843 1 101
2 844 1 101
2 845 1 102
2 846 1 102
2 847 1 103
2 848 1 103
2 849 1 104
2 850 1 104
2 851 1 105
2 852 1 105
2 853 1 106
2 854 1 106
2 855 1 107
2 856 1 107
2 857 1 108
2 858 1 108
2 859 1 109
2 860 1 109
2 861 1 110
2 862 1 110
2 863 1 111
2 864 1 111
2 865 1 112
2 866 1 112
2 867 1 177
2 868 1 177
2 869 1 178
2 870 1 178
2 871 1 179
2 872 1 179
2 873 1 180
2 874 1 180
2 875 1 181
2 876 1 181
2 877 1 182
2 878 1 182
2 879 1 183
2 880 1 183
2 881 1 184
2 882 1 184
2 883 1 185
2 884 1 185
2 885 1 186
2 886 1 186
2 887 1 187
2 888 1 187
2 889 1 188
2 890 1 188
2 891 1 189
2 892 1 189
2 893 1 190
2 894 1 190
2 895 1 191
2 896 1 191
2 897 1 192
2 898 1 192
2 899 1 193
2 900 1 193
2 901 1 194
2 902 1 194
2 903 1 195
2 904 1 195
2 905 1 196
2 906 1 196
2 907 1 197
2 908 1 197
2 909 1 198
2 910 1 198
2 911 1 199
2 912 1 199
2 913 1 200
2 914 1 200
2 915 1 201
2 916 1 201
2 917 1 202
2 918 1 202
2 919 1 203
2 920 1 203
2 921 1 204
2 922 1 204
2 923 1 205
2 924 1 205
2 925 1 206
2 926 1 206
2 927 1 207
2 928 1 207
2 929 1 208
2 930 1 208
2 931 1 209
2 932 1 209
2 933 1 210
2 934 1 210
2 935 1 211
2 936 1 211
2 937 1 212
2 938 1 212
2 939 1 213
2 940 1 213
2 941 1 214
2 942 1 214
2 943 1 215
2 944 1 215
2 945 1 216
2 946 1 216
2 947 1 217
2 948 1 217
2 949 1 218
2 950 1 218
2 951 1 219
2 952 1 219
2 953 1 220
2 954 1 220
2 955 1 221
2 956 1 221
2 957 1 222
2 958 1 222
2 959 1 223
2 960 1 223
2 961 1 224
2 962 1 224
2 963 1 257
2 964 1 257
2 965 1 257
2 966 1 257
2 967 1 258
2 968 1 258
2 969 1 258
2 970 1 258
2 971 1 259
2 972 1 259
2 973 1 259
2 974 1 259
2 975 1 260
2 976 1 260
2 977 1 260
2 978 1 260
2 979 1 261
2 980 1 261
2 981 1 261
2 982 1 261
2 983 1 262
2 984 1 262
2 985 1 262
2 986 1 262
2 987 1 263
2 988 1 263
2 989 1 263
2 990 1 263
2 991 1 264
2 992 1 264
2 993 1 264
2 994 1 264
2 995 1 265
2 996 1 265
2 997 1 266
2 998 1 266
2 999 1 267
2 1000 1 267
2 1001 1 268
2 1002 1 268
2 1003 1 269
2 1004 1 269
2 1005 1 270
2 1006 1 270
2 1007 1 271
2 1008 1 271
2 1009 1 272
2 1010 1 272
2 1011 1 273
2 1012 1 273
2 1013 1 274
2 1014 1 274
2 1015 1 275
2 1016 1 275
2 1017 1 276
2 1018 1 276
2 1019 1 277
2 1020 1 277
2 1021 1 278
2 1022 1 278
2 1023 1 279
2 1024 1 279
2 1025 1 280
2 1026 1 280
2 1027 1 297
2 1028 1 297
2 1029 1 298
2 1030 1 298
2 1031 1 299
2 1032 1 299
2 1033 1 300
2 1034 1 300
2 1035 1 301
2 1036 1 301
2 1037 1 302
2 1038 1 302
2 1039 1 303
2 1040 1 303
2 1041 1 304
2 1042 1 304
2 1043 1 305
2 1044 1 305
2 1045 1 306
2 1046 1 306
2 1047 1 307
2 1048 1 307
2 1049 1 308
2 1050 1 308
2 1051 1 309
2 1052 1 309
2 1053 1 310
2 1054 1 310
2 1055 1 311
2 1056 1 311
2 1057 1 312
2 1058 1 312
2 1059 1 329
2 1060 1 329
2 1061 1 330
2 1062 1 330
2 1063 1 331
2 1064 1 331
2 1065 1 332
2 1066 1 332
2 1067 1 333
2 1068 1 333
2 1069 1 334
2 1070 1 334
2 1071 1 335
2 1072 1 335
2 1073 1 336
2 1074 1 336
2 1075 1 337
2 1076 1 337
2 1077 1 338
2 1078 1 338
2 1079 1 339
2 1080 1 339
2 1081 1 340
2 1082 1 340
2 1083 1 341
2 1084 1 341
2 1085 1 342
2 1086 1 342
2 1087 1 343
2 1088 1 343
2 1089 1 344
2 1090 1 344
2 1091 1 361
2 1092 1 361
2 1093 1 361
2 1094 1 361
2 1095 1 361
2 1096 1 361
2 1097 1 361
2 1098 1 361
2 1099 1 361
2 1100 1 361
2 1101 1 361
2 1102 1 361
2 1103 1 362
2 1104 1 362
2 1105 1 362
2 1106 1 362
2 1107 1 362
2 1108 1 362
2 1109 1 362
2 1110 1 362
2 1111 1 362
2 1112 1 362
2 1113 1 362
2 1114 1 362
2 1115 1 363
2 1116 1 363
2 1117 1 363
2 1118 1 363
2 1119 1 363
2 1120 1 363
2 1121 1 363
2 1122 1 363
2 1123 1 363
2 1124 1 363
2 1125 1 363
2 1126 1 363
2 1127 1 364
2 1128 1 364
2 1129 1 364
2 1130 1 364
2 1131 1 364
2 1132 1 364
2 1133 1 364
2 1134 1 364
2 1135 1 364
2 1136 1 364
2 1137 1 364
2 1138 1 364
2 1139 1 365
2 1140 1 365
2 1141 1 365
2 1142 1 365
2 1143 1 365
2 1144 1 365
2 1145 1 365
2 1146 1 365
2 1147 1 365
2 1148 1 365
2 1149 1 365
2 1150 1 365
2 1151 1 366
2 1152 1 366
2 1153 1 366
2 1154 1 366
2 1155 1 366
2 1156 1 366
2 1157 1 366
2 1158 1 366
2 1159 1 366
2 1160 1 366
2 1161 1 366
2 1162 1 366
2 1163 1 367
2 1164 1 367
2 1165 1 367
2 1166 1 367
2 1167 1 367
2 1168 1 367
2 1169 1 367
2 1170 1 367
2 1171 1 367
2 1172 1 367
2 1173 1 367
2 1174 1 367
2 1175 1 368
2 1176 1 368
2 1177 1 368
2 1178 1 368
2 1179 1 368
2 1180 1 368
2 1181 1 368
2 1182 1 368
2 1183 1 368
2 1184 1 368
2 1185 1 368
2 1186 1 368
2 1187 1 417
2 1188 1 417
2 1189 1 417
2 1190 1 417
2 1191 1 418
2 1192 1 418
2 1193 1 418
2 1194 1 418
2 1195 1 419
2 1196 1 419
2 1197 1 419
2 1198 1 419
2 1199 1 420
2 1200 1 420
2 1201 1 420
2 1202 1 420
2 1203 1 421
2 1204 1 421
2 1205 1 421
2 1206 1 421
2 1207 1 422
2 1208 1 422
2 1209 1 422
2 1210 1 422
2 1211 1 423
2 1212 1 423
2 1213 1 423
2 1214 1 423
2 1215 1 424
2 1216 1 424
2 1217 1 424
2 1218 1 424
2 1219 1 425
2 1220 1 425
2 1221 1 425
2 1222 1 425
2 1223 1 426
2 1224 1 426
2 1225 1 426
2 1226 1 426
2 1227 1 427
2 1228 1 427
2 1229 1 428
2 1230 1 428
2 1231 1 429
2 1232 1 429
2 1233 1 430
2 1234 1 430
2 1235 1 431
2 1236 1 431
2 1237 1 432
2 1238 1 432
2 1239 1 433
2 1240 1 433
2 1241 1 434
2 1242 1 434
2 1243 1 435
2 1244 1 435
2 1245 1 436
2 1246 1 436
2 1247 1 437
2 1248 1 437
2 1249 1 438
2 1250 1 438
2 1251 1 439
2 1252 1 439
2 1253 1 440
2 1254 1 440
2 1255 1 441
2 1256 1 441
2 1257 1 442
2 1258 1 442
2 1259 1 443
2 1260 1 443
2 1261 1 444
2 1262 1 444
2 1263 1 445
2 1264 1 445
2 1265 1 446
2 1266 1 446
2 1267 1 447
2 1268 1 447
2 1269 1 448
2 1270 1 448
2 1271 1 449
2 1272 1 449
2 1273 1 450
2 1274 1 450
2 1275 1 451
2 1276 1 451
2 1277 1 452
2 1278 1 452
2 1279 1 453
2 1280 1 453
2 1281 1 454
2 1282 1 454
2 1283 1 455
2 1284 1 455
2 1285 1 456
2 1286 1 456
2 1287 1 457
2 1288 1 457
2 1289 1 458
2 1290 1 458
2 1291 1 459
2 1292 1 459
2 1293 1 460
2 1294 1 460
2 1295 1 461
2 1296 1 461
2 1297 1 462
2 1298 1 462
2 1299 1 463
2 1300 1 463
2 1301 1 464
2 1302 1 464
2 1303 1 465
2 1304 1 465
2 1305 1 466
2 1306 1 466
2 1307 1 467
2 1308 1 467
2 1309 1 468
2 1310 1 468
2 1311 1 469
2 1312 1 469
2 1313 1 470
2 1314 1 470
2 1315 1 471
2 1316 1 471
2 1317 1 472
2 1318 1 472
2 1319 1 473
2 1320 1 473
2 1321 1 474
2 1322 1 474
2 1323 1 475
2 1324 1 475
2 1325 1 476
2 1326 1 476
2 1327 1 477
2 1328 1 477
2 1329 1 478
2 1330 1 478
2 1331 1 479
2 1332 1 479
2 1333 1 480
2 1334 1 480
2 1335 1 481
2 1336 1 481
2 1337 1 482
2 1338 1 482
2 1339 1 483
2 1340 1 483
2 1341 1 484
2 1342 1 484
2 1343 1 485
2 1344 1 485
2 1345 1 486
2 1346 1 486
2 1347 1 487
2 1348 1 487
2 1349 1 488
2 1350 1 488
2 1351 1 489
2 1352 1 489
2 1353 1 490
2 1354 1 490
