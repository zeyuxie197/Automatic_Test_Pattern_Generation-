1 1 0 1 0
1 2 0 2 0
2 10 1 2
2 11 1 2
1 5 0 1 0
1 6 0 2 0
2 12 1 6
2 13 1 6
1 9 0 1 0
0 14 4 1 2 1 10
0 15 6 2 3 11 12 5
2 19 1 15
2 20 1 15
0 18 5 1 1 13
0 21 4 1 2 18 9
3 22 7 0 2 14 19
3 23 7 0 2 20 21
